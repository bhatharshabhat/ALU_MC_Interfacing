<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>546.421,83.9368,1052.62,-166.268</PageViewport>
<gate>
<ID>1</ID>
<type>AA_AND4</type>
<position>664,17.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>5 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_FULLADDER_1BIT</type>
<position>584.5,-38</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_B_0</ID>9 </input>
<output>
<ID>OUT_0</ID>14 </output>
<input>
<ID>carry_in</ID>10 </input>
<output>
<ID>carry_out</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_FULLADDER_1BIT</type>
<position>567.5,-38</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_B_0</ID>8 </input>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>carry_in</ID>7 </input>
<output>
<ID>carry_out</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>BE_NOR2</type>
<position>821,12.5</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AI_XOR2</type>
<position>566.5,-29</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR2</type>
<position>578.5,-29</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AI_INVERTER_4BIT</type>
<position>658,27.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>1 </input>
<output>
<ID>OUT_0</ID>15 </output>
<output>
<ID>OUT_1</ID>16 </output>
<output>
<ID>OUT_2</ID>23 </output>
<output>
<ID>OUT_3</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>561.5,23.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>561.5,20.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>561.5,17</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>561.5,13.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>555.5,25</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>555.5,21</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>555.5,17.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>555.5,14</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>793.5,-153.5</position>
<output>
<ID>OUT_0</ID>197 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>17</ID>
<type>BE_NOR2</type>
<position>820.5,3.5</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>734,-117.5</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>177 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>561.5,-11</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_OR4</type>
<position>660.5,6.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>5 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>21</ID>
<type>AI_XOR4</type>
<position>662,-4</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>5 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_INVERTER</type>
<position>671.5,12.5</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_INVERTER</type>
<position>674,4</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_INVERTER</type>
<position>673,-8.5</position>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AI_MUX_8x1</type>
<position>691.5,25.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>19 </input>
<input>
<ID>IN_3</ID>11 </input>
<input>
<ID>IN_4</ID>15 </input>
<input>
<ID>IN_5</ID>16 </input>
<input>
<ID>IN_6</ID>23 </input>
<input>
<ID>IN_7</ID>17 </input>
<output>
<ID>OUT</ID>24 </output>
<input>
<ID>SEL_0</ID>13 </input>
<input>
<ID>SEL_1</ID>12 </input>
<input>
<ID>SEL_2</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_MUX_2x1</type>
<position>717.5,24.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>27 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>767.5,24.5</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>BA_DECODER_2x4</type>
<position>775.5,-93</position>
<input>
<ID>IN_0</ID>273 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT_0</ID>151 </output>
<output>
<ID>OUT_1</ID>268 </output>
<output>
<ID>OUT_2</ID>125 </output>
<output>
<ID>OUT_3</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND3</type>
<position>810,11</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>119 </input>
<input>
<ID>IN_2</ID>120 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND3</type>
<position>810,4</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>215 </input>
<input>
<ID>IN_2</ID>120 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>32</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>1050.5,-134.5</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>184 </input>
<input>
<ID>IN_2</ID>185 </input>
<input>
<ID>IN_3</ID>221 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_INVERTER</type>
<position>801.5,11</position>
<input>
<ID>IN_0</ID>215 </input>
<output>
<ID>OUT_0</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>768.5,-113.5</position>
<gparam>LABEL_TEXT A  B</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>608.5,-49</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>608.5,-54</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>768.5,-123.5</position>
<gparam>LABEL_TEXT A = B</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_AND2</type>
<position>608.5,-59</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>768.5,-117.5</position>
<input>
<ID>N_in0</ID>3 </input>
<input>
<ID>N_in1</ID>276 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>608.5,-64</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>769,-134</position>
<gparam>LABEL_TEXT A > B</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AI_XOR2</type>
<position>646.5,-52.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AE_OR4</type>
<position>846,-105</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>143 </input>
<input>
<ID>IN_2</ID>141 </input>
<input>
<ID>IN_3</ID>140 </input>
<output>
<ID>OUT</ID>226 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_AND2</type>
<position>643.5,-57</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AI_MUX_8x1</type>
<position>703.5,-22</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>157 </input>
<input>
<ID>IN_2</ID>157 </input>
<input>
<ID>IN_3</ID>22 </input>
<input>
<ID>IN_4</ID>7 </input>
<input>
<ID>IN_5</ID>14 </input>
<input>
<ID>IN_6</ID>4 </input>
<input>
<ID>IN_7</ID>18 </input>
<output>
<ID>OUT</ID>36 </output>
<input>
<ID>SEL_0</ID>13 </input>
<input>
<ID>SEL_1</ID>12 </input>
<input>
<ID>SEL_2</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>47</ID>
<type>AI_XOR2</type>
<position>655.5,-59.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>769,-128</position>
<input>
<ID>N_in0</ID>40 </input>
<input>
<ID>N_in1</ID>277 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_AND2</type>
<position>656.5,-66.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>767.5,3.5</position>
<input>
<ID>N_in0</ID>37 </input>
<input>
<ID>N_in1</ID>280 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>664.5,-117</position>
<gparam>LABEL_TEXT COMPARATOR</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>GA_LED</type>
<position>769,-138.5</position>
<input>
<ID>N_in0</ID>39 </input>
<input>
<ID>N_in1</ID>278 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>772,-32</position>
<gparam>LABEL_TEXT MUL/ DIV</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_INVERTER</type>
<position>809.5,-2</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>56</ID>
<type>DD_KEYPAD_HEX</type>
<position>563.5,49</position>
<output>
<ID>OUT_0</ID>25 </output>
<output>
<ID>OUT_1</ID>13 </output>
<output>
<ID>OUT_2</ID>12 </output>
<output>
<ID>OUT_3</ID>26 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_AND2</type>
<position>734.5,-128</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>557,30.5</position>
<gparam>LABEL_TEXT INPUTS</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_AND3</type>
<position>835.5,12.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>121 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_AND2</type>
<position>735,-138.5</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>179 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_OR4</type>
<position>907.5,-105.5</position>
<input>
<ID>IN_0</ID>191 </input>
<input>
<ID>IN_1</ID>187 </input>
<input>
<ID>IN_2</ID>169 </input>
<input>
<ID>IN_3</ID>163 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_OR4</type>
<position>975,-105</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>204 </input>
<input>
<ID>IN_2</ID>201 </input>
<input>
<ID>IN_3</ID>195 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>64</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>577.5,33</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>5 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>766.5,32</position>
<gparam>LABEL_TEXT Output</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AE_OR4</type>
<position>1043.5,-105</position>
<input>
<ID>IN_0</ID>217 </input>
<input>
<ID>IN_1</ID>214 </input>
<input>
<ID>IN_2</ID>211 </input>
<input>
<ID>IN_3</ID>207 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>765,7.5</position>
<gparam>LABEL_TEXT Int. C/ B</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>578,3</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>6 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>560,-4.5</position>
<gparam>LABEL_TEXT Key A/ S</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>846,-116</position>
<input>
<ID>N_in2</ID>181 </input>
<input>
<ID>N_in3</ID>226 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>576.5,76.5</position>
<gparam>LABEL_TEXT ALPHANUMERIC OPCODES</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>GA_LED</type>
<position>907.5,-116</position>
<input>
<ID>N_in2</ID>184 </input>
<input>
<ID>N_in3</ID>224 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>584.5,67</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>12 </input>
<input>
<ID>IN_3</ID>26 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>975,-116</position>
<input>
<ID>N_in2</ID>185 </input>
<input>
<ID>N_in3</ID>230 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>BE_NOR2</type>
<position>821,-30.5</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>BE_NOR2</type>
<position>821,-41</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_AND3</type>
<position>809.5,-32</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>127 </input>
<output>
<ID>OUT</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_AND3</type>
<position>812,-40</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>276 </input>
<input>
<ID>IN_2</ID>127 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>98</ID>
<type>GA_LED</type>
<position>1043.5,-115.5</position>
<input>
<ID>N_in3</ID>221 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_INVERTER</type>
<position>801.5,-32</position>
<input>
<ID>IN_0</ID>276 </input>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>770,-60</position>
<gparam>LABEL_TEXT DECODER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AA_INVERTER</type>
<position>812.5,-46</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_AND3</type>
<position>836,-30.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>128 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>797.5,-162</position>
<gparam>LABEL_TEXT READ / WRITE</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_AND3</type>
<position>663.5,-71.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>49 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_INVERTER</type>
<position>656.5,-73.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_OR2</type>
<position>659,-78.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_AND3</type>
<position>670.5,-81.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>1 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND3</type>
<position>668,-87.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>51 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_INVERTER</type>
<position>656,-90.5</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR3</type>
<position>714.5,-80</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>54 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_LABEL</type>
<position>805.5,-156</position>
<gparam>LABEL_TEXT ________</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND3</type>
<position>668.5,-95</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>56 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_INVERTER</type>
<position>646,-96.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>123</ID>
<type>BE_NOR2</type>
<position>883,12</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>137 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>BE_NOR2</type>
<position>883,3</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>618.5,-30</position>
<gparam>LABEL_TEXT ADDER/ SUB</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>631,-65.5</position>
<gparam>LABEL_TEXT MULTIPLIER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_AND3</type>
<position>872.5,10.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>133 </input>
<input>
<ID>IN_2</ID>269 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_LABEL</type>
<position>604,-78.5</position>
<gparam>LABEL_TEXT DIVIDER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_AND3</type>
<position>872.5,3.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>245 </input>
<input>
<ID>IN_2</ID>269 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_LABEL</type>
<position>1039.5,-141.5</position>
<gparam>LABEL_TEXT OUTPUT </gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_INVERTER</type>
<position>861.5,10.5</position>
<input>
<ID>IN_0</ID>245 </input>
<output>
<ID>OUT_0</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_INVERTER</type>
<position>872.5,-2</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>269 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND3</type>
<position>897.5,13</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>136 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>151</ID>
<type>BE_NOR2</type>
<position>884,-29</position>
<input>
<ID>IN_0</ID>138 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>152</ID>
<type>BE_NOR2</type>
<position>884,-39</position>
<input>
<ID>IN_0</ID>145 </input>
<input>
<ID>IN_1</ID>139 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_AND3</type>
<position>872.5,-31.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>142 </input>
<input>
<ID>IN_2</ID>144 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>156</ID>
<type>AA_AND3</type>
<position>872.5,-38.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>277 </input>
<input>
<ID>IN_2</ID>144 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>158</ID>
<type>AA_INVERTER</type>
<position>862,-31.5</position>
<input>
<ID>IN_0</ID>277 </input>
<output>
<ID>OUT_0</ID>142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_INVERTER</type>
<position>873,-44</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>162</ID>
<type>AA_AND3</type>
<position>898,-28.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>145 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>166</ID>
<type>BE_NOR2</type>
<position>815.5,51.5</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>162 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>BE_NOR2</type>
<position>816,43</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND3</type>
<position>807.5,50.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>158 </input>
<input>
<ID>IN_2</ID>160 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_AND3</type>
<position>807.5,43</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>134 </input>
<input>
<ID>IN_2</ID>160 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_INVERTER</type>
<position>799.5,50.5</position>
<input>
<ID>IN_0</ID>134 </input>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_INVERTER</type>
<position>806.5,37</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_AND3</type>
<position>835,51.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>161 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>180</ID>
<type>FF_GND</type>
<position>919,-4.5</position>
<output>
<ID>OUT_0</ID>271 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_AND3</type>
<position>609.5,-100.5</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_2</ID>2 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>184</ID>
<type>BE_NOR2</type>
<position>883,49</position>
<input>
<ID>IN_0</ID>164 </input>
<input>
<ID>IN_1</ID>275 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_AND2</type>
<position>609.5,-107.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>186</ID>
<type>BE_NOR2</type>
<position>883,40</position>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>165 </input>
<output>
<ID>OUT</ID>275 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_AND3</type>
<position>609.5,-114</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>2 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_AND3</type>
<position>872.5,47.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>186 </input>
<input>
<ID>IN_2</ID>188 </input>
<output>
<ID>OUT</ID>164 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>189</ID>
<type>AE_OR3</type>
<position>637.5,-118.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>86 </input>
<input>
<ID>IN_2</ID>87 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_AND3</type>
<position>872.5,40.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>149 </input>
<input>
<ID>IN_2</ID>188 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_INVERTER</type>
<position>590,-98.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_INVERTER</type>
<position>862.5,47.5</position>
<input>
<ID>IN_0</ID>149 </input>
<output>
<ID>OUT_0</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>193</ID>
<type>AA_INVERTER</type>
<position>593.5,-102.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_INVERTER</type>
<position>872,35</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>195</ID>
<type>AA_INVERTER</type>
<position>591.5,-106.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_AND3</type>
<position>897.5,49</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>189 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_INVERTER</type>
<position>591.5,-112</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>198</ID>
<type>FF_GND</type>
<position>986.5,-4.5</position>
<output>
<ID>OUT_0</ID>270 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>199</ID>
<type>BE_NOR2</type>
<position>823.5,-74.5</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>274 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>BE_NOR2</type>
<position>823.5,-82.5</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>274 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>AO_XNOR2</type>
<position>609.5,-121</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_AND3</type>
<position>810,-75.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>196 </input>
<input>
<ID>IN_2</ID>198 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>203</ID>
<type>AO_XNOR2</type>
<position>609.5,-126</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_AND3</type>
<position>810,-82.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>198 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_AND2</type>
<position>637,-129</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_INVERTER</type>
<position>801,-75.5</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_AND3</type>
<position>609,-134</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>97 </input>
<input>
<ID>IN_2</ID>98 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_INVERTER</type>
<position>810,-88</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_AND3</type>
<position>609,-141</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>1 </input>
<input>
<ID>IN_2</ID>99 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_AND3</type>
<position>836.5,-74.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>199 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_AND2</type>
<position>609,-147</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>AE_OR3</type>
<position>638,-139.5</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>110 </input>
<input>
<ID>IN_2</ID>111 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>214</ID>
<type>BE_NOR2</type>
<position>885.5,-75.5</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>210 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>BE_NOR2</type>
<position>885.5,-84.5</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>203 </input>
<output>
<ID>OUT</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_AND3</type>
<position>874.5,-77</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>206 </input>
<input>
<ID>IN_2</ID>208 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_INVERTER</type>
<position>591,-134</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_AND3</type>
<position>874.5,-84</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>22 </input>
<input>
<ID>IN_2</ID>208 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>219</ID>
<type>AA_INVERTER</type>
<position>597,-136</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_INVERTER</type>
<position>862.5,-77</position>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_INVERTER</type>
<position>596,-143</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_INVERTER</type>
<position>874,-89.5</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>208 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>223</ID>
<type>AA_INVERTER</type>
<position>591,-148</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_AND3</type>
<position>898.5,-74.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>209 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>225</ID>
<type>FF_GND</type>
<position>985,-48.5</position>
<output>
<ID>OUT_0</ID>279 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>226</ID>
<type>BE_NOR2</type>
<position>949.5,50</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>220 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>BE_NOR2</type>
<position>949.5,41</position>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>213 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_AND3</type>
<position>937.5,48.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>216 </input>
<input>
<ID>IN_2</ID>218 </input>
<output>
<ID>OUT</ID>212 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_AND3</type>
<position>937.5,41.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>148 </input>
<input>
<ID>IN_2</ID>218 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_INVERTER</type>
<position>926.5,48.5</position>
<input>
<ID>IN_0</ID>148 </input>
<output>
<ID>OUT_0</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>231</ID>
<type>AA_INVERTER</type>
<position>936.5,36</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>218 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_AND3</type>
<position>964.5,50</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>219 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>234</ID>
<type>BE_NOR2</type>
<position>951.5,11</position>
<input>
<ID>IN_0</ID>222 </input>
<input>
<ID>IN_1</ID>229 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>235</ID>
<type>BE_NOR2</type>
<position>951.5,1.5</position>
<input>
<ID>IN_0</ID>228 </input>
<input>
<ID>IN_1</ID>223 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND3</type>
<position>939.5,8.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>225 </input>
<input>
<ID>IN_2</ID>227 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>237</ID>
<type>AA_AND3</type>
<position>939.5,1.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>271 </input>
<input>
<ID>IN_2</ID>227 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>238</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>774,-40.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>149 </input>
<input>
<ID>IN_2</ID>148 </input>
<input>
<ID>IN_3</ID>152 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_INVERTER</type>
<position>926.5,8.5</position>
<input>
<ID>IN_0</ID>271 </input>
<output>
<ID>OUT_0</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_AND2</type>
<position>732.5,-34</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>AA_INVERTER</type>
<position>939,-4</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>227 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>242</ID>
<type>AA_AND2</type>
<position>732.5,-39</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_AND3</type>
<position>964,11</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>228 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>244</ID>
<type>AA_AND2</type>
<position>732.5,-44</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>245</ID>
<type>FF_GND</type>
<position>988,-81.5</position>
<output>
<ID>OUT_0</ID>281 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_AND2</type>
<position>732.5,-49</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>180 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>247</ID>
<type>BE_NOR2</type>
<position>951,-26.5</position>
<input>
<ID>IN_0</ID>231 </input>
<input>
<ID>IN_1</ID>236 </input>
<output>
<ID>OUT</ID>235 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>BE_NOR2</type>
<position>951,-37</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>232 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>249</ID>
<type>AA_AND3</type>
<position>939.5,-29.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>233 </input>
<input>
<ID>IN_2</ID>234 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_AND3</type>
<position>939.5,-36.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>278 </input>
<input>
<ID>IN_2</ID>234 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_INVERTER</type>
<position>924.5,-29.5</position>
<input>
<ID>IN_0</ID>278 </input>
<output>
<ID>OUT_0</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_INVERTER</type>
<position>939,-42</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>234 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_AND3</type>
<position>964.5,-26</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>235 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>255</ID>
<type>BE_NOR2</type>
<position>950,-70.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>241 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_INVERTER</type>
<position>717,-13.5</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>153 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>257</ID>
<type>BE_NOR2</type>
<position>950,-80</position>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_AND3</type>
<position>939,-73</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>239 </input>
<input>
<ID>IN_2</ID>240 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>259</ID>
<type>AA_AND3</type>
<position>939,-80</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>280 </input>
<input>
<ID>IN_2</ID>240 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>260</ID>
<type>AA_INVERTER</type>
<position>721.5,-14.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_INVERTER</type>
<position>923.5,-73</position>
<input>
<ID>IN_0</ID>280 </input>
<output>
<ID>OUT_0</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_INVERTER</type>
<position>725.5,-10.5</position>
<input>
<ID>IN_0</ID>25 </input>
<output>
<ID>OUT_0</ID>155 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_INVERTER</type>
<position>938.5,-85.5</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>240 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_AND4</type>
<position>720,-29.5</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>12 </input>
<input>
<ID>IN_3</ID>153 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_AND3</type>
<position>965.5,-70.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>241 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>195 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>266</ID>
<type>FF_GND</type>
<position>698.5,-36</position>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>267</ID>
<type>AA_TOGGLE</type>
<position>756.5,-153.5</position>
<output>
<ID>OUT_0</ID>273 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>268</ID>
<type>BE_NOR2</type>
<position>1017.5,53.5</position>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_1</ID>249 </input>
<output>
<ID>OUT</ID>248 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>269</ID>
<type>BE_NOR2</type>
<position>1017.5,42.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>249 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>270</ID>
<type>AA_AND3</type>
<position>1006.5,50</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>246 </input>
<input>
<ID>IN_2</ID>247 </input>
<output>
<ID>OUT</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_AND3</type>
<position>1006.5,42.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>152 </input>
<input>
<ID>IN_2</ID>247 </input>
<output>
<ID>OUT</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_INVERTER</type>
<position>992.5,50</position>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT_0</ID>246 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_INVERTER</type>
<position>1006,37</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>247 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>274</ID>
<type>AA_AND3</type>
<position>1034.5,54</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>248 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_INVERTER</type>
<position>724,-71.5</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>277</ID>
<type>BE_NOR2</type>
<position>1016.5,10</position>
<input>
<ID>IN_0</ID>250 </input>
<input>
<ID>IN_1</ID>255 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_INVERTER</type>
<position>728.5,-71.5</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>167 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>279</ID>
<type>BE_NOR2</type>
<position>1016.5,2</position>
<input>
<ID>IN_0</ID>254 </input>
<input>
<ID>IN_1</ID>251 </input>
<output>
<ID>OUT</ID>255 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_INVERTER</type>
<position>733,-72</position>
<input>
<ID>IN_0</ID>25 </input>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>281</ID>
<type>AA_AND3</type>
<position>1004.5,8.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>252 </input>
<input>
<ID>IN_2</ID>253 </input>
<output>
<ID>OUT</ID>250 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>282</ID>
<type>AA_AND4</type>
<position>727,-86.5</position>
<input>
<ID>IN_0</ID>168 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>167 </input>
<input>
<ID>IN_3</ID>166 </input>
<output>
<ID>OUT</ID>170 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>283</ID>
<type>AA_AND3</type>
<position>1004.5,1.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>270 </input>
<input>
<ID>IN_2</ID>253 </input>
<output>
<ID>OUT</ID>251 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>284</ID>
<type>AA_INVERTER</type>
<position>993,8.5</position>
<input>
<ID>IN_0</ID>270 </input>
<output>
<ID>OUT_0</ID>252 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>285</ID>
<type>AA_INVERTER</type>
<position>1004,-4</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>253 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>286</ID>
<type>AA_AND2</type>
<position>735,-91</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>287</ID>
<type>AA_AND3</type>
<position>1034.5,10</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>254 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_AND2</type>
<position>735,-97.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>289</ID>
<type>AA_TOGGLE</type>
<position>750.5,-153.5</position>
<output>
<ID>OUT_0</ID>272 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>290</ID>
<type>AA_INVERTER</type>
<position>685,-102</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>172 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>291</ID>
<type>BE_NOR2</type>
<position>1015,-29</position>
<input>
<ID>IN_0</ID>256 </input>
<input>
<ID>IN_1</ID>261 </input>
<output>
<ID>OUT</ID>260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>292</ID>
<type>AA_INVERTER</type>
<position>689.5,-101</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>173 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>293</ID>
<type>BE_NOR2</type>
<position>1015,-40</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>257 </input>
<output>
<ID>OUT</ID>261 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>294</ID>
<type>AA_INVERTER</type>
<position>693.5,-103</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>174 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>295</ID>
<type>AA_AND3</type>
<position>1004,-31.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>258 </input>
<input>
<ID>IN_2</ID>259 </input>
<output>
<ID>OUT</ID>256 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>296</ID>
<type>AA_INVERTER</type>
<position>698,-101.5</position>
<input>
<ID>IN_0</ID>25 </input>
<output>
<ID>OUT_0</ID>175 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>297</ID>
<type>AA_AND3</type>
<position>1004,-38.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>279 </input>
<input>
<ID>IN_2</ID>259 </input>
<output>
<ID>OUT</ID>257 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_AND4</type>
<position>691.5,-115</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>174 </input>
<input>
<ID>IN_2</ID>173 </input>
<input>
<ID>IN_3</ID>172 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>299</ID>
<type>AA_INVERTER</type>
<position>992,-31.5</position>
<input>
<ID>IN_0</ID>279 </input>
<output>
<ID>OUT_0</ID>258 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>300</ID>
<type>AE_OR2</type>
<position>747.5,-57.5</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>301</ID>
<type>AA_INVERTER</type>
<position>1003.5,-44.5</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>259 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>302</ID>
<type>AE_OR2</type>
<position>747.5,-64</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>245 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>AA_AND3</type>
<position>1033.5,-28.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>260 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>305</ID>
<type>BE_NOR2</type>
<position>1015,-70</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>267 </input>
<output>
<ID>OUT</ID>266 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>BE_NOR2</type>
<position>1015,-79.5</position>
<input>
<ID>IN_0</ID>266 </input>
<input>
<ID>IN_1</ID>263 </input>
<output>
<ID>OUT</ID>267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>AA_AND3</type>
<position>1004.5,-71.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>264 </input>
<input>
<ID>IN_2</ID>265 </input>
<output>
<ID>OUT</ID>262 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>308</ID>
<type>AA_AND3</type>
<position>1004.5,-78.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>281 </input>
<input>
<ID>IN_2</ID>265 </input>
<output>
<ID>OUT</ID>263 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>309</ID>
<type>AA_INVERTER</type>
<position>992.5,-71.5</position>
<input>
<ID>IN_0</ID>281 </input>
<output>
<ID>OUT_0</ID>264 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>310</ID>
<type>AA_INVERTER</type>
<position>1004,-84.5</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>265 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>311</ID>
<type>AA_AND3</type>
<position>1034,-70</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>266 </input>
<input>
<ID>IN_2</ID>197 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_LABEL</type>
<position>760,-159.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>313</ID>
<type>AA_LABEL</type>
<position>747,-159.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>315</ID>
<type>AA_LABEL</type>
<position>832.5,-115.5</position>
<gparam>LABEL_TEXT OP0</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>316</ID>
<type>AA_LABEL</type>
<position>893.5,-115</position>
<gparam>LABEL_TEXT OP1</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>317</ID>
<type>AA_LABEL</type>
<position>961.5,-116</position>
<gparam>LABEL_TEXT OP2</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>318</ID>
<type>AA_LABEL</type>
<position>1030.5,-116</position>
<gparam>LABEL_TEXT OP3</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>324</ID>
<type>AA_LABEL</type>
<position>821.5,69</position>
<gparam>LABEL_TEXT 4x4 RAM</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>326</ID>
<type>AA_LABEL</type>
<position>643.5,65.5</position>
<gparam>LABEL_TEXT ALU</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>624,-12.5,624,23.5</points>
<intersection>-12.5 28</intersection>
<intersection>-1 26</intersection>
<intersection>9.5 14</intersection>
<intersection>21.5 4</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>563.5,23.5,656,23.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>573 54</intersection>
<intersection>624 0</intersection>
<intersection>656 50</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>624,21.5,659.5,21.5</points>
<intersection>624 0</intersection>
<intersection>659.5 51</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>624,9.5,657.5,9.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>624 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>624,-1,659,-1</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>624 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>601,-12.5,624,-12.5</points>
<intersection>601 30</intersection>
<intersection>624 0</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>601,-48,601,-12.5</points>
<intersection>-48 31</intersection>
<intersection>-35 32</intersection>
<intersection>-12.5 28</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>593.5,-48,605.5,-48</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>593.5 33</intersection>
<intersection>601 30</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>585.5,-35,601,-35</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>601 30</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>593.5,-58,593.5,-48</points>
<intersection>-58 34</intersection>
<intersection>-48 31</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>572.5,-58,605.5,-58</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>572.5 36</intersection>
<intersection>593.5 33</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>572.5,-69.5,572.5,-58</points>
<intersection>-69.5 37</intersection>
<intersection>-58 34</intersection></vsegment>
<hsegment>
<ID>37</ID>
<points>561,-69.5,660.5,-69.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>561 38</intersection>
<intersection>572.5 36</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>561,-83.5,561,-69.5</points>
<intersection>-83.5 39</intersection>
<intersection>-69.5 37</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>561,-83.5,667.5,-83.5</points>
<connection>
<GID>115</GID>
<name>IN_2</name></connection>
<intersection>561 38</intersection>
<intersection>567.5 40</intersection></hsegment>
<vsegment>
<ID>40</ID>
<points>567.5,-102.5,567.5,-83.5</points>
<intersection>-102.5 41</intersection>
<intersection>-83.5 39</intersection></vsegment>
<hsegment>
<ID>41</ID>
<points>559,-102.5,590.5,-102.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>559 42</intersection>
<intersection>567.5 40</intersection></hsegment>
<vsegment>
<ID>42</ID>
<points>559,-141,559,-102.5</points>
<intersection>-141 49</intersection>
<intersection>-132 47</intersection>
<intersection>-125 45</intersection>
<intersection>-112 43</intersection>
<intersection>-102.5 41</intersection></vsegment>
<hsegment>
<ID>43</ID>
<points>559,-112,588.5,-112</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>559 42</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>559,-125,606.5,-125</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>559 42</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>559,-132,606,-132</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>559 42</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>559,-141,606,-141</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>559 42</intersection></hsegment>
<vsegment>
<ID>50</ID>
<points>656,23.5,656,29</points>
<connection>
<GID>7</GID>
<name>IN_3</name></connection>
<intersection>23.5 1</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>659.5,20.5,659.5,21.5</points>
<intersection>20.5 52</intersection>
<intersection>21.5 4</intersection></vsegment>
<hsegment>
<ID>52</ID>
<points>659.5,20.5,661,20.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>659.5 51</intersection></hsegment>
<vsegment>
<ID>54</ID>
<points>573,23.5,573,32</points>
<intersection>23.5 1</intersection>
<intersection>32 55</intersection></vsegment>
<hsegment>
<ID>55</ID>
<points>573,32,574.5,32</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>573 54</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>627,-19,627,28</points>
<intersection>-19 26</intersection>
<intersection>-3 23</intersection>
<intersection>7.5 14</intersection>
<intersection>20.5 2</intersection>
<intersection>28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>627,28,656,28</points>
<connection>
<GID>7</GID>
<name>IN_2</name></connection>
<intersection>627 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>563.5,20.5,654,20.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>567.5 60</intersection>
<intersection>627 0</intersection>
<intersection>654 56</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>627,7.5,657.5,7.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>627 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>627,-3,659,-3</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>627 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>577.5,-19,627,-19</points>
<intersection>577.5 27</intersection>
<intersection>598 33</intersection>
<intersection>627 0</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>577.5,-26,577.5,-19</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-19 26</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>598,-50,598,-19</points>
<intersection>-50 34</intersection>
<intersection>-19 26</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>598,-50,605.5,-50</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>598 33</intersection>
<intersection>601 35</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>601,-55,601,-50</points>
<intersection>-55 36</intersection>
<intersection>-50 34</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>562.5,-55,605.5,-55</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>562.5 38</intersection>
<intersection>601 35</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>562.5,-71.5,562.5,-55</points>
<intersection>-71.5 39</intersection>
<intersection>-55 36</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>562.5,-71.5,660.5,-71.5</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>562.5 38</intersection>
<intersection>636.5 40</intersection></hsegment>
<vsegment>
<ID>40</ID>
<points>636.5,-77.5,636.5,-71.5</points>
<intersection>-77.5 41</intersection>
<intersection>-71.5 39</intersection></vsegment>
<hsegment>
<ID>41</ID>
<points>615.5,-77.5,656,-77.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>615.5 42</intersection>
<intersection>636.5 40</intersection></hsegment>
<vsegment>
<ID>42</ID>
<points>615.5,-90.5,615.5,-77.5</points>
<intersection>-90.5 43</intersection>
<intersection>-77.5 41</intersection></vsegment>
<hsegment>
<ID>43</ID>
<points>563,-90.5,653,-90.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>563 44</intersection>
<intersection>615.5 42</intersection></hsegment>
<vsegment>
<ID>44</ID>
<points>563,-95,563,-90.5</points>
<intersection>-95 45</intersection>
<intersection>-90.5 43</intersection></vsegment>
<hsegment>
<ID>45</ID>
<points>563,-95,665.5,-95</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>563 44</intersection>
<intersection>573.5 46</intersection></hsegment>
<vsegment>
<ID>46</ID>
<points>573.5,-104.5,573.5,-95</points>
<intersection>-104.5 47</intersection>
<intersection>-95 45</intersection></vsegment>
<hsegment>
<ID>47</ID>
<points>564.5,-104.5,597.5,-104.5</points>
<intersection>564.5 48</intersection>
<intersection>573.5 46</intersection>
<intersection>597.5 57</intersection></hsegment>
<vsegment>
<ID>48</ID>
<points>564.5,-143,564.5,-104.5</points>
<intersection>-143 55</intersection>
<intersection>-136 53</intersection>
<intersection>-127 51</intersection>
<intersection>-116 49</intersection>
<intersection>-104.5 47</intersection></vsegment>
<hsegment>
<ID>49</ID>
<points>564.5,-116,606.5,-116</points>
<connection>
<GID>187</GID>
<name>IN_2</name></connection>
<intersection>564.5 48</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>564.5,-127,606.5,-127</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>564.5 48</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>564.5,-136,594,-136</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>564.5 48</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>564.5,-143,593,-143</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>564.5 48</intersection></hsegment>
<vsegment>
<ID>56</ID>
<points>654,18.5,654,20.5</points>
<intersection>18.5 59</intersection>
<intersection>20.5 2</intersection></vsegment>
<vsegment>
<ID>57</ID>
<points>597.5,-104.5,597.5,-102.5</points>
<intersection>-104.5 47</intersection>
<intersection>-102.5 58</intersection></vsegment>
<hsegment>
<ID>58</ID>
<points>597.5,-102.5,606.5,-102.5</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>597.5 57</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>654,18.5,661,18.5</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>654 56</intersection></hsegment>
<vsegment>
<ID>60</ID>
<points>567.5,2,567.5,20.5</points>
<intersection>2 61</intersection>
<intersection>20.5 2</intersection></vsegment>
<hsegment>
<ID>61</ID>
<points>567.5,2,575,2</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>567.5 60</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>737,-117.5,767.5,-117.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>688,-19.5,688,-8.5</points>
<intersection>-19.5 3</intersection>
<intersection>-8.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>688,-19.5,700.5,-19.5</points>
<connection>
<GID>46</GID>
<name>IN_6</name></connection>
<intersection>688 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>676,-8.5,688,-8.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>688 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>630.5,-16.5,630.5,27</points>
<intersection>-16.5 28</intersection>
<intersection>-5 26</intersection>
<intersection>5.5 18</intersection>
<intersection>17 15</intersection>
<intersection>27 22</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>563.5,17,661,17</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>571.5 54</intersection>
<intersection>630.5 0</intersection>
<intersection>661 35</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>630.5,5.5,657.5,5.5</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>630.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>630.5,27,656,27</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>630.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>630.5,-5,659,-5</points>
<connection>
<GID>21</GID>
<name>IN_2</name></connection>
<intersection>630.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>559,-16.5,630.5,-16.5</points>
<intersection>559 30</intersection>
<intersection>630.5 0</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>559,-98.5,559,-16.5</points>
<intersection>-98.5 44</intersection>
<intersection>-85.5 40</intersection>
<intersection>-81.5 38</intersection>
<intersection>-53 31</intersection>
<intersection>-35 32</intersection>
<intersection>-16.5 28</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>559,-53,605.5,-53</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>559 30</intersection>
<intersection>582 33</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>559,-35,568.5,-35</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>559 30</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>582,-63,582,-53</points>
<intersection>-63 34</intersection>
<intersection>-53 31</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>566,-63,605.5,-63</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>566 37</intersection>
<intersection>582 33</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>661,16.5,661,17</points>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>17 15</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>566,-81.5,566,-63</points>
<intersection>-81.5 38</intersection>
<intersection>-63 34</intersection></vsegment>
<hsegment>
<ID>38</ID>
<points>559,-81.5,667.5,-81.5</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>559 30</intersection>
<intersection>566 37</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>559,-85.5,665,-85.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>559 30</intersection>
<intersection>614 41</intersection></hsegment>
<vsegment>
<ID>41</ID>
<points>614,-93,614,-85.5</points>
<intersection>-93 42</intersection>
<intersection>-85.5 40</intersection></vsegment>
<hsegment>
<ID>42</ID>
<points>614,-93,665.5,-93</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>614 41</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>559,-98.5,587,-98.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>559 30</intersection>
<intersection>583.5 45</intersection></hsegment>
<vsegment>
<ID>45</ID>
<points>583.5,-106.5,583.5,-98.5</points>
<intersection>-106.5 46</intersection>
<intersection>-98.5 44</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>567,-106.5,588.5,-106.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>567 47</intersection>
<intersection>583.5 45</intersection></hsegment>
<vsegment>
<ID>47</ID>
<points>567,-146,567,-106.5</points>
<intersection>-146 52</intersection>
<intersection>-139 50</intersection>
<intersection>-120 48</intersection>
<intersection>-106.5 46</intersection></vsegment>
<hsegment>
<ID>48</ID>
<points>567,-120,606.5,-120</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>567 47</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>567,-139,606,-139</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>567 47</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>567,-146,606,-146</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>567 47</intersection></hsegment>
<vsegment>
<ID>54</ID>
<points>571.5,17,571.5,33</points>
<intersection>17 15</intersection>
<intersection>33 55</intersection></vsegment>
<hsegment>
<ID>55</ID>
<points>571.5,33,574.5,33</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>571.5 54</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>634.5,-7,634.5,26</points>
<intersection>-7 4</intersection>
<intersection>3.5 7</intersection>
<intersection>14.5 6</intersection>
<intersection>26 24</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>620.5,-7,659,-7</points>
<connection>
<GID>21</GID>
<name>IN_3</name></connection>
<intersection>620.5 12</intersection>
<intersection>634.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>634.5,14.5,661,14.5</points>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>634.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>634.5,3.5,657.5,3.5</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<intersection>634.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>620.5,-16.5,620.5,13.5</points>
<intersection>-16.5 21</intersection>
<intersection>-7 4</intersection>
<intersection>13.5 27</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>565.5,-16.5,620.5,-16.5</points>
<intersection>565.5 22</intersection>
<intersection>600 28</intersection>
<intersection>620.5 12</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>565.5,-26,565.5,-16.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>-16.5 21</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>634.5,26,656,26</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>634.5 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>563.5,13.5,620.5,13.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>569 49</intersection>
<intersection>620.5 12</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>600,-65,600,-16.5</points>
<intersection>-65 30</intersection>
<intersection>-60 29</intersection>
<intersection>-16.5 21</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>600,-60,605.5,-60</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>600 28</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>588,-65,605.5,-65</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>588 31</intersection>
<intersection>600 28</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>588,-73.5,588,-65</points>
<intersection>-73.5 32</intersection>
<intersection>-65 30</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>588,-73.5,653.5,-73.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>588 31</intersection>
<intersection>648 33</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>648,-79.5,648,-73.5</points>
<intersection>-79.5 34</intersection>
<intersection>-73.5 32</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>624.5,-79.5,656,-79.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>624.5 35</intersection>
<intersection>648 33</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>624.5,-87.5,624.5,-79.5</points>
<intersection>-87.5 36</intersection>
<intersection>-79.5 34</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>561,-87.5,665,-87.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>561 37</intersection>
<intersection>624.5 35</intersection></hsegment>
<vsegment>
<ID>37</ID>
<points>561,-148,561,-87.5</points>
<intersection>-148 48</intersection>
<intersection>-134 46</intersection>
<intersection>-122 44</intersection>
<intersection>-114 42</intersection>
<intersection>-108.5 40</intersection>
<intersection>-96.5 38</intersection>
<intersection>-87.5 36</intersection></vsegment>
<hsegment>
<ID>38</ID>
<points>561,-96.5,643,-96.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>561 37</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>561,-108.5,606.5,-108.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>561 37</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>561,-114,606.5,-114</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>561 37</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>561,-122,606.5,-122</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>561 37</intersection>
<intersection>584.5 45</intersection></hsegment>
<vsegment>
<ID>45</ID>
<points>584.5,-134,584.5,-122</points>
<intersection>-134 46</intersection>
<intersection>-122 44</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>561,-134,588,-134</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>561 37</intersection>
<intersection>584.5 45</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>561,-148,588,-148</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>561 37</intersection></hsegment>
<vsegment>
<ID>49</ID>
<points>569,3,569,13.5</points>
<intersection>3 50</intersection>
<intersection>13.5 27</intersection></vsegment>
<hsegment>
<ID>50</ID>
<points>569,3,575,3</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>569 49</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>571.5,-43,693.5,-43</points>
<intersection>571.5 14</intersection>
<intersection>580.5 13</intersection>
<intersection>693.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>693.5,-43,693.5,-21.5</points>
<intersection>-43 6</intersection>
<intersection>-21.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>693.5,-21.5,700.5,-21.5</points>
<connection>
<GID>46</GID>
<name>IN_4</name></connection>
<intersection>693.5 9</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>580.5,-43,580.5,-38</points>
<connection>
<GID>2</GID>
<name>carry_out</name></connection>
<intersection>-43 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>571.5,-43,571.5,-38</points>
<connection>
<GID>3</GID>
<name>carry_in</name></connection>
<intersection>-43 6</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>566.5,-35,566.5,-32</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<connection>
<GID>3</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583.5,-35,583.5,-32</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<intersection>-32 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>578.5,-32,583.5,-32</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>583.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593.5,-38,593.5,-11</points>
<intersection>-38 3</intersection>
<intersection>-24.5 4</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>563.5,-11,593.5,-11</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>567.5 2</intersection>
<intersection>593.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>567.5,-26,567.5,-11</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>588.5,-38,593.5,-38</points>
<connection>
<GID>2</GID>
<name>carry_in</name></connection>
<intersection>593.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>579.5,-24.5,593.5,-24.5</points>
<intersection>579.5 5</intersection>
<intersection>593.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>579.5,-26,579.5,-24.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-24.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>667,17.5,677,17.5</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<intersection>667 4</intersection>
<intersection>677 13</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>667,12.5,667,17.5</points>
<intersection>12.5 5</intersection>
<intersection>17.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>667,12.5,668.5,12.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>667 4</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>677,17.5,677,25</points>
<intersection>17.5 1</intersection>
<intersection>25 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>677,25,688.5,25</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>677 13</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>703.5,-16.5,703.5,50</points>
<connection>
<GID>46</GID>
<name>SEL_1</name></connection>
<intersection>-7 15</intersection>
<intersection>50 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>568.5,50,703.5,50</points>
<connection>
<GID>56</GID>
<name>OUT_2</name></connection>
<intersection>571.5 25</intersection>
<intersection>691.5 11</intersection>
<intersection>703.5 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>691.5,31,691.5,50</points>
<connection>
<GID>25</GID>
<name>SEL_1</name></connection>
<intersection>50 6</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>703.5,-7,708,-7</points>
<intersection>703.5 0</intersection>
<intersection>708 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>708,-38,708,-7</points>
<intersection>-38 17</intersection>
<intersection>-26.5 21</intersection>
<intersection>-7 15</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>689.5,-38,708,-38</points>
<intersection>689.5 18</intersection>
<intersection>708 16</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>689.5,-98,689.5,-38</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>-61 19</intersection>
<intersection>-38 17</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>689.5,-61,728.5,-61</points>
<intersection>689.5 18</intersection>
<intersection>728.5 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>728.5,-68.5,728.5,-61</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>-61 19</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>708,-26.5,719,-26.5</points>
<connection>
<GID>264</GID>
<name>IN_2</name></connection>
<intersection>708 16</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>571.5,50,571.5,68</points>
<intersection>50 6</intersection>
<intersection>68 26</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>571.5,68,581.5,68</points>
<connection>
<GID>80</GID>
<name>IN_2</name></connection>
<intersection>571.5 25</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>706,-16.5,706,48</points>
<intersection>-16.5 33</intersection>
<intersection>-4 20</intersection>
<intersection>48 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>568.5,48,706,48</points>
<connection>
<GID>56</GID>
<name>OUT_1</name></connection>
<intersection>573 36</intersection>
<intersection>692.5 16</intersection>
<intersection>706 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>692.5,31,692.5,48</points>
<connection>
<GID>25</GID>
<name>SEL_0</name></connection>
<intersection>48 15</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>682.5,-4,706,-4</points>
<intersection>682.5 21</intersection>
<intersection>706 0</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>682.5,-54,682.5,-4</points>
<intersection>-54 22</intersection>
<intersection>-11.5 23</intersection>
<intersection>-4 20</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>682.5,-54,731,-54</points>
<intersection>682.5 21</intersection>
<intersection>731 24</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>682.5,-11.5,721.5,-11.5</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>682.5 21</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>731,-54,731,-52</points>
<intersection>-54 22</intersection>
<intersection>-52 25</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>693.5,-52,731,-52</points>
<intersection>693.5 26</intersection>
<intersection>731 24</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>693.5,-100,693.5,-52</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>-83.5 29</intersection>
<intersection>-52 25</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>693.5,-83.5,728,-83.5</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<intersection>693.5 26</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>704.5,-16.5,706,-16.5</points>
<connection>
<GID>46</GID>
<name>SEL_0</name></connection>
<intersection>706 0</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>573,48,573,67</points>
<intersection>48 15</intersection>
<intersection>67 37</intersection></vsegment>
<hsegment>
<ID>37</ID>
<points>573,67,581.5,67</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>573 36</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584.5,-41,584.5,-20.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>556,-20.5,700.5,-20.5</points>
<connection>
<GID>46</GID>
<name>IN_5</name></connection>
<intersection>556 2</intersection>
<intersection>584.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>556,-75.5,556,-20.5</points>
<intersection>-75.5 3</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>556,-75.5,798,-75.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>556 2</intersection>
<intersection>796.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>796.5,-82.5,796.5,-75.5</points>
<intersection>-82.5 5</intersection>
<intersection>-75.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>796.5,-82.5,807,-82.5</points>
<connection>
<GID>204</GID>
<name>IN_1</name></connection>
<intersection>796.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>660,26,688.5,26</points>
<connection>
<GID>25</GID>
<name>IN_4</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>660,27,688.5,27</points>
<connection>
<GID>25</GID>
<name>IN_5</name></connection>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>660,29,688.5,29</points>
<connection>
<GID>25</GID>
<name>IN_7</name></connection>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>666,-4,670,-4</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>670 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>670,-18.5,670,-4</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-18.5 11</intersection>
<intersection>-4 7</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>670,-18.5,700.5,-18.5</points>
<connection>
<GID>46</GID>
<name>IN_7</name></connection>
<intersection>670 9</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>679,24,688.5,24</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>679 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>679,12.5,679,24</points>
<intersection>12.5 5</intersection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>674.5,12.5,679,12.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>679 4</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>664.5,6.5,681.5,6.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>664.5 3</intersection>
<intersection>681.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>664.5,4,664.5,6.5</points>
<intersection>4 4</intersection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>664.5,4,671,4</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>664.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>681.5,6.5,681.5,23</points>
<intersection>6.5 1</intersection>
<intersection>23 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>681.5,23,688.5,23</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>681.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>684.5,4,684.5,22</points>
<intersection>4 3</intersection>
<intersection>22 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>677,4,684.5,4</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>684.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>684.5,22,688.5,22</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>684.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>569.5,-41,569.5,-22.5</points>
<intersection>-41 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>569.5,-22.5,856,-22.5</points>
<connection>
<GID>46</GID>
<name>IN_3</name></connection>
<intersection>569.5 0</intersection>
<intersection>856 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>567.5,-41,569.5,-41</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>569.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>856,-84,856,-22.5</points>
<intersection>-84 6</intersection>
<intersection>-77 4</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>856,-77,859.5,-77</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>856 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>856,-84,871.5,-84</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>856 3</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>660,28,688.5,28</points>
<connection>
<GID>25</GID>
<name>IN_6</name></connection>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>694.5,25.5,715.5,25.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<connection>
<GID>25</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>709.5,29.5,709.5,46</points>
<intersection>29.5 1</intersection>
<intersection>46 16</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>709.5,29.5,736.5,29.5</points>
<intersection>709.5 0</intersection>
<intersection>717.5 3</intersection>
<intersection>736.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>736.5,-2,736.5,29.5</points>
<intersection>-2 6</intersection>
<intersection>29.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>717.5,27,717.5,29.5</points>
<connection>
<GID>26</GID>
<name>SEL_0</name></connection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>680.5,-2,736.5,-2</points>
<intersection>680.5 7</intersection>
<intersection>736.5 2</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>680.5,-58,680.5,-2</points>
<intersection>-58 8</intersection>
<intersection>-6 9</intersection>
<intersection>-2 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>680.5,-58,707.5,-58</points>
<intersection>680.5 7</intersection>
<intersection>707.5 10</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>680.5,-6,725.5,-6</points>
<intersection>680.5 7</intersection>
<intersection>725.5 11</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>707.5,-98.5,707.5,-58</points>
<intersection>-98.5 12</intersection>
<intersection>-67.5 13</intersection>
<intersection>-58 8</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>725.5,-7.5,725.5,-6</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>-6 9</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>698,-98.5,707.5,-98.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>707.5 10</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>707.5,-67.5,733,-67.5</points>
<intersection>707.5 10</intersection>
<intersection>733 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>733,-69,733,-67.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>-67.5 13</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>568.5,46,709.5,46</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>574.5 20</intersection>
<intersection>709.5 0</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>574.5,46,574.5,66</points>
<intersection>46 16</intersection>
<intersection>66 21</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>574.5,66,581.5,66</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>574.5 20</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>701,-16.5,701,52</points>
<intersection>-16.5 31</intersection>
<intersection>-10.5 15</intersection>
<intersection>52 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>568.5,52,701,52</points>
<connection>
<GID>56</GID>
<name>OUT_3</name></connection>
<intersection>570 35</intersection>
<intersection>690.5 13</intersection>
<intersection>701 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>690.5,31,690.5,52</points>
<connection>
<GID>25</GID>
<name>SEL_2</name></connection>
<intersection>52 6</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>677.5,-10.5,717,-10.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>677.5 22</intersection>
<intersection>701 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>677.5,-97.5,677.5,-10.5</points>
<intersection>-97.5 25</intersection>
<intersection>-65 23</intersection>
<intersection>-10.5 15</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>677.5,-65,724,-65</points>
<intersection>677.5 22</intersection>
<intersection>724 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>724,-68.5,724,-65</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>-65 23</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>677.5,-97.5,685,-97.5</points>
<intersection>677.5 22</intersection>
<intersection>685 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>685,-99,685,-97.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>-97.5 25</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>701,-16.5,702.5,-16.5</points>
<connection>
<GID>46</GID>
<name>SEL_2</name></connection>
<intersection>701 0</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>570,52,570,69</points>
<intersection>52 6</intersection>
<intersection>69 36</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>570,69,581.5,69</points>
<connection>
<GID>80</GID>
<name>IN_3</name></connection>
<intersection>570 35</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>719.5,24.5,766.5,24.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>27</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>623,-54,623,-51.5</points>
<intersection>-54 2</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>623,-51.5,643.5,-51.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>623 0</intersection>
<intersection>635.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>611.5,-54,623,-54</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>623 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>635.5,-56,635.5,-51.5</points>
<intersection>-56 4</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>635.5,-56,640.5,-56</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>635.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>624.5,-59,624.5,-53.5</points>
<intersection>-59 2</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>624.5,-53.5,643.5,-53.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>624.5 0</intersection>
<intersection>631.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>611.5,-59,624.5,-59</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>624.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>631.5,-58,631.5,-53.5</points>
<intersection>-58 4</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>631.5,-58,640.5,-58</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>631.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>647.5,-58.5,647.5,-57</points>
<intersection>-58.5 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>647.5,-58.5,652.5,-58.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>647.5 0</intersection>
<intersection>649.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>646.5,-57,647.5,-57</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>647.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>649.5,-65.5,649.5,-58.5</points>
<intersection>-65.5 4</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>649.5,-65.5,653.5,-65.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>649.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>630,-64,630,-60.5</points>
<intersection>-64 2</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>630,-60.5,652.5,-60.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>630 0</intersection>
<intersection>646.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>611.5,-64,630,-64</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>630 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>646.5,-67.5,646.5,-60.5</points>
<intersection>-67.5 4</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>646.5,-67.5,653.5,-67.5</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>646.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>673,-56,673,-49</points>
<intersection>-56 1</intersection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>673,-56,729,-56</points>
<intersection>673 0</intersection>
<intersection>729 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>611.5,-49,673,-49</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<intersection>673 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>729,-56,729,-50</points>
<intersection>-56 1</intersection>
<intersection>-50 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>729,-50,729.5,-50</points>
<connection>
<GID>246</GID>
<name>IN_1</name></connection>
<intersection>729 5</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>691.5,-63,691.5,-52.5</points>
<intersection>-63 1</intersection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>691.5,-63,717,-63</points>
<intersection>691.5 0</intersection>
<intersection>717 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>649.5,-52.5,691.5,-52.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>691.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>717,-63,717,-45</points>
<intersection>-63 1</intersection>
<intersection>-45 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>717,-45,729.5,-45</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>717 5</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>698,-69,698,-59.5</points>
<intersection>-69 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>698,-69,715.5,-69</points>
<intersection>698 0</intersection>
<intersection>715.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>658.5,-59.5,698,-59.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>698 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>715.5,-69,715.5,-40</points>
<intersection>-69 1</intersection>
<intersection>-40 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>715.5,-40,729.5,-40</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>715.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>659.5,-66.5,714,-66.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>714 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>714,-66.5,714,-35</points>
<intersection>-66.5 1</intersection>
<intersection>-35 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>714,-35,729.5,-35</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>714 7</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>710,-22,710,23.5</points>
<intersection>-22 3</intersection>
<intersection>23.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>706.5,-22,710,-22</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>710 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>710,23.5,715.5,23.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>710 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>563.5,-46,712,-46</points>
<intersection>563.5 4</intersection>
<intersection>712 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>712,-46,712,3.5</points>
<intersection>-46 1</intersection>
<intersection>3.5 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>563.5,-46,563.5,-38</points>
<connection>
<GID>3</GID>
<name>carry_out</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>712,3.5,766.5,3.5</points>
<connection>
<GID>50</GID>
<name>N_in0</name></connection>
<intersection>712 3</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>738,-138.5,768,-138.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<connection>
<GID>53</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>737.5,-128,768,-128</points>
<connection>
<GID>57</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>659.5,-73.5,660.5,-73.5</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<connection>
<GID>112</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>662,-78.5,665,-78.5</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>665 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>665,-79.5,665,-78.5</points>
<intersection>-79.5 3</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>665,-79.5,667.5,-79.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>665 2</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>660.5,-89.5,665,-89.5</points>
<connection>
<GID>116</GID>
<name>IN_2</name></connection>
<intersection>660.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>660.5,-90.5,660.5,-89.5</points>
<intersection>-90.5 6</intersection>
<intersection>-89.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>659,-90.5,660.5,-90.5</points>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<intersection>660.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673.5,-81.5,708.5,-81.5</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>708.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>708.5,-81.5,708.5,-80</points>
<intersection>-81.5 1</intersection>
<intersection>-80 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>708.5,-80,711.5,-80</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>708.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>692.5,-78,692.5,-71.5</points>
<intersection>-78 1</intersection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>692.5,-78,711.5,-78</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>692.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>666.5,-71.5,692.5,-71.5</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>692.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>671,-87.5,708.5,-87.5</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>708.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>708.5,-87.5,708.5,-82</points>
<intersection>-87.5 1</intersection>
<intersection>-82 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>708.5,-82,711.5,-82</points>
<connection>
<GID>118</GID>
<name>IN_2</name></connection>
<intersection>708.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>720,-103,720,-80</points>
<intersection>-103 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>720,-103,731,-103</points>
<intersection>720 0</intersection>
<intersection>731 9</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>717.5,-80,720,-80</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>720 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>731,-103,731,-98.5</points>
<intersection>-103 1</intersection>
<intersection>-98.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>731,-98.5,732,-98.5</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<intersection>731 9</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649,-96.5,665.5,-96.5</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>665.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>665.5,-97,665.5,-96.5</points>
<connection>
<GID>120</GID>
<name>IN_2</name></connection>
<intersection>-96.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>715.5,-104.5,715.5,-95</points>
<intersection>-104.5 1</intersection>
<intersection>-95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>715.5,-104.5,730,-104.5</points>
<intersection>715.5 0</intersection>
<intersection>730 9</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>671.5,-95,715.5,-95</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>715.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>730,-104.5,730,-92</points>
<intersection>-104.5 1</intersection>
<intersection>-92 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>730,-92,732,-92</points>
<connection>
<GID>286</GID>
<name>IN_1</name></connection>
<intersection>730 9</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>631.5,-116.5,631.5,-100.5</points>
<intersection>-116.5 1</intersection>
<intersection>-100.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>631.5,-116.5,634.5,-116.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>631.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>612.5,-100.5,631.5,-100.5</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<intersection>631.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612.5,-107.5,629.5,-107.5</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>629.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>629.5,-118.5,629.5,-107.5</points>
<intersection>-118.5 3</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>629.5,-118.5,634.5,-118.5</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<intersection>629.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>622.5,-120.5,622.5,-114</points>
<intersection>-120.5 2</intersection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>612.5,-114,622.5,-114</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<intersection>622.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>622.5,-120.5,634.5,-120.5</points>
<connection>
<GID>189</GID>
<name>IN_2</name></connection>
<intersection>622.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593,-98.5,606.5,-98.5</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<connection>
<GID>183</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>597,-100.5,606.5,-100.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>597 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>597,-102.5,597,-100.5</points>
<intersection>-102.5 9</intersection>
<intersection>-100.5 0</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>596.5,-102.5,597,-102.5</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<intersection>597 8</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>594.5,-106.5,606.5,-106.5</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<connection>
<GID>185</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>594.5,-112,606.5,-112</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>594,-134,606,-134</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600,-136,606,-136</points>
<connection>
<GID>207</GID>
<name>IN_2</name></connection>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>599,-143,606,-143</points>
<connection>
<GID>209</GID>
<name>IN_2</name></connection>
<connection>
<GID>221</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>594,-148,606,-148</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>621,-128,621,-121</points>
<intersection>-128 1</intersection>
<intersection>-121 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>621,-128,634,-128</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>621 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>612.5,-121,621,-121</points>
<connection>
<GID>201</GID>
<name>OUT</name></connection>
<intersection>621 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>614,-130,634,-130</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>614 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>614,-130,614,-126</points>
<intersection>-130 1</intersection>
<intersection>-126 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>612.5,-126,614,-126</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>614 3</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612,-137.5,635,-137.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>612 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>612,-137.5,612,-134</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<intersection>-137.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>623,-141,623,-139.5</points>
<intersection>-141 2</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>623,-139.5,635,-139.5</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>623 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>612,-141,623,-141</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<intersection>623 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>624,-147,624,-141.5</points>
<intersection>-147 2</intersection>
<intersection>-141.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>624,-141.5,635,-141.5</points>
<connection>
<GID>213</GID>
<name>IN_2</name></connection>
<intersection>624 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>612,-147,624,-147</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>624 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>813,13.5,818,13.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>813 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>813,11,813,13.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>813,2.5,817.5,2.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>813 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>813,2.5,813,4</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>2.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>804.5,11,807,11</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<connection>
<GID>29</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>801,-2,801,9</points>
<intersection>-2 1</intersection>
<intersection>2 2</intersection>
<intersection>9 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>801,-2,806.5,-2</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>801 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>801,2,807,2</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<intersection>801 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>801,9,807,9</points>
<connection>
<GID>29</GID>
<name>IN_2</name></connection>
<intersection>801 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>824,12.5,832.5,12.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>824.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>824.5,7,824.5,12.5</points>
<intersection>7 4</intersection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>814.5,7,824.5,7</points>
<intersection>814.5 5</intersection>
<intersection>824.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>814.5,4.5,814.5,7</points>
<intersection>4.5 9</intersection>
<intersection>7 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>814.5,4.5,817.5,4.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>814.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>823.5,3.5,826,3.5</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>826 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>826,3.5,826,9</points>
<intersection>3.5 1</intersection>
<intersection>9 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>815,9,826,9</points>
<intersection>815 5</intersection>
<intersection>826 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>815,9,815,11.5</points>
<intersection>9 4</intersection>
<intersection>11.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>815,11.5,818,11.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>815 5</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>815,-32,815,-29.5</points>
<intersection>-32 8</intersection>
<intersection>-29.5 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>812.5,-32,815,-32</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>815 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>815,-29.5,818,-29.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>815 7</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>815,-42,818,-42</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<intersection>815 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>815,-42,815,-40</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>805,-38,805,-20.5</points>
<intersection>-38 1</intersection>
<intersection>-30 56</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>805,-38,809,-38</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>805 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>786.5,-20.5,1022,-20.5</points>
<intersection>786.5 57</intersection>
<intersection>805 0</intersection>
<intersection>827 5</intersection>
<intersection>867 14</intersection>
<intersection>890.5 19</intersection>
<intersection>931 28</intersection>
<intersection>957.5 33</intersection>
<intersection>998 42</intersection>
<intersection>1022 47</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>827,-28.5,827,-20.5</points>
<intersection>-28.5 7</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>827,-28.5,833,-28.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>827 5</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>867,-39.5,867,-16</points>
<intersection>-39.5 15</intersection>
<intersection>-20.5 2</intersection>
<intersection>-16 26</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>867,-39.5,1001,-39.5</points>
<intersection>867 14</intersection>
<intersection>869.5 63</intersection>
<intersection>998 42</intersection>
<intersection>1001 64</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>890.5,-26.5,890.5,-20.5</points>
<intersection>-26.5 21</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>890.5,-26.5,895,-26.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>890.5 19</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>867,-16,1001,-16</points>
<intersection>867 14</intersection>
<intersection>869.5 60</intersection>
<intersection>957.5 33</intersection>
<intersection>961.5 62</intersection>
<intersection>998 42</intersection>
<intersection>1001 61</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>931,-34.5,931,-20.5</points>
<intersection>-34.5 29</intersection>
<intersection>-27.5 40</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>931,-34.5,936.5,-34.5</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>931 28</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>957.5,-20.5,957.5,-16</points>
<intersection>-20.5 2</intersection>
<intersection>-16 26</intersection></vsegment>
<hsegment>
<ID>40</ID>
<points>931,-27.5,936.5,-27.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>931 28</intersection></hsegment>
<vsegment>
<ID>42</ID>
<points>998,-39.5,998,-16</points>
<intersection>-39.5 15</intersection>
<intersection>-20.5 2</intersection>
<intersection>-16 26</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>1022,-26.5,1022,-20.5</points>
<intersection>-26.5 49</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>49</ID>
<points>1022,-26.5,1030.5,-26.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>1022 47</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>805,-30,806.5,-30</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>805 0</intersection></hsegment>
<vsegment>
<ID>57</ID>
<points>786.5,-92.5,786.5,-20.5</points>
<intersection>-92.5 58</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>58</ID>
<points>778.5,-92.5,786.5,-92.5</points>
<connection>
<GID>28</GID>
<name>OUT_2</name></connection>
<intersection>786.5 57</intersection></hsegment>
<vsegment>
<ID>60</ID>
<points>869.5,-29.5,869.5,-16</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>-16 26</intersection></vsegment>
<vsegment>
<ID>61</ID>
<points>1001,-29.5,1001,-16</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>-16 26</intersection></vsegment>
<vsegment>
<ID>62</ID>
<points>961.5,-24,961.5,-16</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>-16 26</intersection></vsegment>
<vsegment>
<ID>63</ID>
<points>869.5,-39.5,869.5,-36.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-39.5 15</intersection></vsegment>
<vsegment>
<ID>64</ID>
<points>1001,-39.5,1001,-36.5</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>-39.5 15</intersection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>804.5,-32,806.5,-32</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<connection>
<GID>94</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>803.5,-46,803.5,-34</points>
<intersection>-46 1</intersection>
<intersection>-42 2</intersection>
<intersection>-34 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>803.5,-46,809.5,-46</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>803.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>803.5,-42,809,-42</points>
<connection>
<GID>96</GID>
<name>IN_2</name></connection>
<intersection>803.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>803.5,-34,806.5,-34</points>
<connection>
<GID>94</GID>
<name>IN_2</name></connection>
<intersection>803.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>824,-30.5,833,-30.5</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>825.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>825.5,-36.5,825.5,-30.5</points>
<intersection>-36.5 4</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>816.5,-36.5,825.5,-36.5</points>
<intersection>816.5 5</intersection>
<intersection>825.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>816.5,-40,816.5,-36.5</points>
<intersection>-40 9</intersection>
<intersection>-36.5 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>816.5,-40,818,-40</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>816.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>824,-41,827,-41</points>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>827 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>827,-41,827,-33.5</points>
<intersection>-41 1</intersection>
<intersection>-33.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>816.5,-33.5,827,-33.5</points>
<intersection>816.5 5</intersection>
<intersection>827 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>816.5,-33.5,816.5,-31.5</points>
<intersection>-33.5 4</intersection>
<intersection>-31.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>816.5,-31.5,818,-31.5</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>816.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>875.5,13,880,13</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>875.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>875.5,10.5,875.5,13</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<intersection>13 1</intersection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>875.5,2,880,2</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>875.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>875.5,2,875.5,3.5</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>2 1</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>864.5,10.5,869.5,10.5</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<connection>
<GID>128</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>760.5,-57.5,760.5,-41.5</points>
<intersection>-57.5 2</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>749,-41.5,771,-41.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>749 3</intersection>
<intersection>760.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>750.5,-57.5,760.5,-57.5</points>
<connection>
<GID>300</GID>
<name>OUT</name></connection>
<intersection>760.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>749,-41.5,749,72</points>
<intersection>-41.5 1</intersection>
<intersection>72 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>749,72,792,72</points>
<intersection>749 3</intersection>
<intersection>792 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>792,43,792,72</points>
<intersection>43 8</intersection>
<intersection>50.5 6</intersection>
<intersection>72 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>792,50.5,796.5,50.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>792 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>792,43,804.5,43</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<intersection>792 5</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>886,13,894.5,13</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>886 22</intersection>
<intersection>889 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>889,7,889,13</points>
<intersection>7 4</intersection>
<intersection>13 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>877,7,889,7</points>
<intersection>877 5</intersection>
<intersection>889 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>877,4,877,7</points>
<intersection>4 9</intersection>
<intersection>7 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>877,4,880,4</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>877 5</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>886,12,886,13</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>13 1</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>886,3,887,3</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<intersection>887 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>887,3,887,9</points>
<intersection>3 1</intersection>
<intersection>9 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>877,9,887,9</points>
<intersection>877 5</intersection>
<intersection>887 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>877,9,877,11</points>
<intersection>9 4</intersection>
<intersection>11 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>877,11,880,11</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>877 5</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>875.5,-28,881,-28</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>875.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>875.5,-31.5,875.5,-28</points>
<connection>
<GID>154</GID>
<name>OUT</name></connection>
<intersection>-28 1</intersection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>875.5,-40,881,-40</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>875.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>875.5,-40,875.5,-38.5</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<intersection>-40 1</intersection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>843,-102,843,-74.5</points>
<connection>
<GID>44</GID>
<name>IN_3</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>839.5,-74.5,843,-74.5</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<intersection>843 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>845,-102,845,-30.5</points>
<connection>
<GID>44</GID>
<name>IN_2</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>839,-30.5,845,-30.5</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<intersection>845 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>865,-31.5,869.5,-31.5</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<connection>
<GID>154</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>847,-102,847,12.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>838.5,12.5,847,12.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>847 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>863,-44,863,-33.5</points>
<intersection>-44 1</intersection>
<intersection>-40.5 2</intersection>
<intersection>-33.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>863,-44,870,-44</points>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection>
<intersection>863 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>863,-40.5,869.5,-40.5</points>
<connection>
<GID>156</GID>
<name>IN_2</name></connection>
<intersection>863 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>863,-33.5,869.5,-33.5</points>
<connection>
<GID>154</GID>
<name>IN_2</name></connection>
<intersection>863 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>887,-28.5,895,-28.5</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>887 10</intersection>
<intersection>889 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>889,-34.5,889,-28.5</points>
<intersection>-34.5 4</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>877,-34.5,889,-34.5</points>
<intersection>877 5</intersection>
<intersection>889 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>877,-38,877,-34.5</points>
<intersection>-38 9</intersection>
<intersection>-34.5 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>877,-38,881,-38</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>877 5</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>887,-29,887,-28.5</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<intersection>-28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>887,-39,888,-39</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<intersection>888 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>888,-39,888,-33</points>
<intersection>-39 1</intersection>
<intersection>-33 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>877,-33,888,-33</points>
<intersection>877 5</intersection>
<intersection>888 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>877,-33,877,-30</points>
<intersection>-33 4</intersection>
<intersection>-30 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>877,-30,881,-30</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<intersection>877 5</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>810.5,52.5,812.5,52.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>810.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>810.5,50.5,810.5,52.5</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<intersection>52.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>735.5,-39.5,771,-39.5</points>
<connection>
<GID>238</GID>
<name>IN_2</name></connection>
<intersection>735.5 3</intersection>
<intersection>744 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>735.5,-39.5,735.5,-39</points>
<connection>
<GID>242</GID>
<name>OUT</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>744,-39.5,744,77</points>
<intersection>-39.5 1</intersection>
<intersection>77 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>744,77,920,77</points>
<intersection>744 4</intersection>
<intersection>920 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>920,41.5,920,77</points>
<intersection>41.5 10</intersection>
<intersection>48.5 7</intersection>
<intersection>77 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>920,48.5,923.5,48.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>920 6</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>920,41.5,934.5,41.5</points>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<intersection>920 6</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>752,-64,752,-40.5</points>
<intersection>-64 2</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>746.5,-40.5,771,-40.5</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<intersection>746.5 3</intersection>
<intersection>752 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>750.5,-64,752,-64</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<intersection>752 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>746.5,-40.5,746.5,74.5</points>
<intersection>-40.5 1</intersection>
<intersection>74.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>746.5,74.5,856,74.5</points>
<intersection>746.5 3</intersection>
<intersection>856 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>856,40.5,856,74.5</points>
<intersection>40.5 8</intersection>
<intersection>47.5 6</intersection>
<intersection>74.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>856,47.5,859.5,47.5</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>856 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>856,40.5,869.5,40.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>856 5</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>810.5,42,813,42</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>810.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>810.5,42,810.5,43</points>
<connection>
<GID>172</GID>
<name>OUT</name></connection>
<intersection>42 1</intersection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>788.5,-94.5,788.5,60.5</points>
<intersection>-94.5 13</intersection>
<intersection>45 1</intersection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>788.5,45,804.5,45</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>788.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>788.5,60.5,1024.5,60.5</points>
<intersection>788.5 0</intersection>
<intersection>803.5 56</intersection>
<intersection>820.5 5</intersection>
<intersection>866.5 15</intersection>
<intersection>887 20</intersection>
<intersection>931.5 29</intersection>
<intersection>956 34</intersection>
<intersection>998 43</intersection>
<intersection>1024.5 48</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>820.5,53.5,820.5,60.5</points>
<intersection>53.5 7</intersection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>820.5,53.5,832,53.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>820.5 5</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>778.5,-94.5,788.5,-94.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>788.5 0</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>866.5,42.5,866.5,60.5</points>
<intersection>42.5 16</intersection>
<intersection>49.5 27</intersection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>866.5,42.5,869.5,42.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>866.5 15</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>887,51,887,60.5</points>
<intersection>51 22</intersection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>887,51,894.5,51</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>887 20</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>866.5,49.5,869.5,49.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>866.5 15</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>931.5,43.5,931.5,60.5</points>
<intersection>43.5 30</intersection>
<intersection>50.5 41</intersection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>931.5,43.5,934.5,43.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>931.5 29</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>956,52,956,60.5</points>
<intersection>52 36</intersection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>956,52,1003.5,52</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>956 34</intersection>
<intersection>998 43</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>931.5,50.5,934.5,50.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>931.5 29</intersection></hsegment>
<vsegment>
<ID>43</ID>
<points>998,44.5,998,60.5</points>
<intersection>44.5 44</intersection>
<intersection>52 36</intersection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>44</ID>
<points>998,44.5,1003.5,44.5</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>998 43</intersection></hsegment>
<vsegment>
<ID>48</ID>
<points>1024.5,56,1024.5,60.5</points>
<intersection>56 50</intersection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>50</ID>
<points>1024.5,56,1031.5,56</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>1024.5 48</intersection></hsegment>
<vsegment>
<ID>56</ID>
<points>803.5,52.5,803.5,60.5</points>
<intersection>52.5 57</intersection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>57</ID>
<points>803.5,52.5,804.5,52.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>803.5 56</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>741.5,-38.5,741.5,79.5</points>
<intersection>-38.5 1</intersection>
<intersection>-34 2</intersection>
<intersection>79.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>741.5,-38.5,771,-38.5</points>
<connection>
<GID>238</GID>
<name>IN_3</name></connection>
<intersection>741.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>735.5,-34,741.5,-34</points>
<connection>
<GID>240</GID>
<name>OUT</name></connection>
<intersection>741.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>741.5,79.5,985.5,79.5</points>
<intersection>741.5 0</intersection>
<intersection>985.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>985.5,42.5,985.5,79.5</points>
<intersection>42.5 6</intersection>
<intersection>50 7</intersection>
<intersection>79.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>985.5,42.5,1003.5,42.5</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<intersection>985.5 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>985.5,50,989.5,50</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>985.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>717,-26.5,717,-16.5</points>
<connection>
<GID>264</GID>
<name>IN_3</name></connection>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>721,-26.5,721,-19</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>721,-19,721.5,-19</points>
<intersection>721 0</intersection>
<intersection>721.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>721.5,-19,721.5,-17.5</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<intersection>-19 2</intersection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>723,-26.5,723,-20.5</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>725.5,-20.5,725.5,-13.5</points>
<connection>
<GID>262</GID>
<name>OUT_0</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>723,-20.5,725.5,-20.5</points>
<intersection>723 0</intersection>
<intersection>725.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>720,-48,720,-32.5</points>
<connection>
<GID>264</GID>
<name>OUT</name></connection>
<intersection>-48 7</intersection>
<intersection>-43 5</intersection>
<intersection>-38 3</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>720,-33,729.5,-33</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>720 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>720,-38,729.5,-38</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>720 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>720,-43,729.5,-43</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>720 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>720,-48,729.5,-48</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>720 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>698.5,-35,698.5,-23.5</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 1</intersection>
<intersection>-24.5 5</intersection>
<intersection>-23.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>698.5,-25.5,700.5,-25.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>698.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>698.5,-24.5,700.5,-24.5</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>698.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>698.5,-23.5,700.5,-23.5</points>
<connection>
<GID>46</GID>
<name>IN_2</name></connection>
<intersection>698.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>802.5,50.5,804.5,50.5</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>849,-102,849,51.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>838,51.5,849,51.5</points>
<connection>
<GID>178</GID>
<name>OUT</name></connection>
<intersection>849 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>800,37,800,48.5</points>
<intersection>37 1</intersection>
<intersection>41 2</intersection>
<intersection>48.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>800,37,803.5,37</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>800 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>800,41,804.5,41</points>
<connection>
<GID>172</GID>
<name>IN_2</name></connection>
<intersection>800 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>800,48.5,804.5,48.5</points>
<connection>
<GID>170</GID>
<name>IN_2</name></connection>
<intersection>800 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>818.5,51.5,832,51.5</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>822.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>822.5,46,822.5,51.5</points>
<intersection>46 4</intersection>
<intersection>51.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>811,46,822.5,46</points>
<intersection>811 5</intersection>
<intersection>822.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>811,44,811,46</points>
<intersection>44 9</intersection>
<intersection>46 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>811,44,813,44</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>811 5</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>819,43,821,43</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<intersection>821 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>821,43,821,47</points>
<intersection>43 1</intersection>
<intersection>47 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>811,47,821,47</points>
<intersection>811 5</intersection>
<intersection>821 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>811,47,811,50.5</points>
<intersection>47 4</intersection>
<intersection>50.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>811,50.5,812.5,50.5</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>811 5</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>904.5,-102.5,904.5,-74.5</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>901.5,-74.5,904.5,-74.5</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<intersection>904.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>875.5,50,880,50</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>875.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>875.5,47.5,875.5,50</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>50 1</intersection></vsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>875.5,39,880,39</points>
<connection>
<GID>186</GID>
<name>IN_1</name></connection>
<intersection>875.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>875.5,39,875.5,40.5</points>
<connection>
<GID>190</GID>
<name>OUT</name></connection>
<intersection>39 1</intersection></vsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>724,-83.5,724,-74.5</points>
<connection>
<GID>282</GID>
<name>IN_3</name></connection>
<connection>
<GID>276</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>726,-83.5,726,-77</points>
<connection>
<GID>282</GID>
<name>IN_2</name></connection>
<intersection>-77 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>728.5,-77,728.5,-74.5</points>
<connection>
<GID>278</GID>
<name>OUT_0</name></connection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>726,-77,728.5,-77</points>
<intersection>726 0</intersection>
<intersection>728.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>733,-78.5,733,-75</points>
<connection>
<GID>280</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>730,-78.5,733,-78.5</points>
<intersection>730 4</intersection>
<intersection>733 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>730,-83.5,730,-78.5</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>-78.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>906.5,-102.5,906.5,-28.5</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>901,-28.5,906.5,-28.5</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>906.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>727,-96.5,727,-89.5</points>
<connection>
<GID>282</GID>
<name>OUT</name></connection>
<intersection>-96.5 3</intersection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>727,-90,732,-90</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>727 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>727,-96.5,732,-96.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>727 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>688.5,-112,688.5,-105</points>
<connection>
<GID>298</GID>
<name>IN_3</name></connection>
<intersection>-105 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>685,-105,688.5,-105</points>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection>
<intersection>688.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>689.5,-104,690.5,-104</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<intersection>690.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>690.5,-112,690.5,-104</points>
<connection>
<GID>298</GID>
<name>IN_2</name></connection>
<intersection>-104 5</intersection></vsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>692.5,-112,692.5,-106</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>-106 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>692.5,-106,693.5,-106</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>692.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>694.5,-112,694.5,-104.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>-104.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>694.5,-104.5,698,-104.5</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<intersection>694.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>691.5,-119,691.5,-118</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>691.5,-119,698.5,-119</points>
<intersection>691.5 0</intersection>
<intersection>698.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>698.5,-119,698.5,-116.5</points>
<intersection>-119 1</intersection>
<intersection>-116.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>698.5,-116.5,731,-116.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>698.5 2</intersection>
<intersection>713.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>713.5,-137.5,713.5,-116.5</points>
<intersection>-137.5 7</intersection>
<intersection>-127 5</intersection>
<intersection>-116.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>713.5,-127,731.5,-127</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>713.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>713.5,-137.5,732,-137.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>713.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>644,-122,716,-122</points>
<intersection>644 4</intersection>
<intersection>716 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>716,-122,716,-118.5</points>
<intersection>-122 1</intersection>
<intersection>-118.5 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>644,-122,644,-118.5</points>
<intersection>-122 1</intersection>
<intersection>-118.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>716,-118.5,731,-118.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>716 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>640.5,-118.5,644,-118.5</points>
<connection>
<GID>189</GID>
<name>OUT</name></connection>
<intersection>644 4</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>640,-129,731.5,-129</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<connection>
<GID>205</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>641,-139.5,732,-139.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<connection>
<GID>213</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>741.5,-56.5,741.5,-49</points>
<intersection>-56.5 2</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>735.5,-49,741.5,-49</points>
<connection>
<GID>246</GID>
<name>OUT</name></connection>
<intersection>741.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>741.5,-56.5,744.5,-56.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>741.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>846,-135.5,846,-117</points>
<connection>
<GID>70</GID>
<name>N_in2</name></connection>
<intersection>-135.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>846,-135.5,1047.5,-135.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>846 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>742.5,-63,742.5,-44</points>
<intersection>-63 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>735.5,-44,742.5,-44</points>
<connection>
<GID>244</GID>
<name>OUT</name></connection>
<intersection>742.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>742.5,-63,744.5,-63</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>742.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>907.5,-134.5,907.5,-117</points>
<connection>
<GID>76</GID>
<name>N_in2</name></connection>
<intersection>-134.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>907.5,-134.5,1047.5,-134.5</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>907.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>975,-133.5,975,-117</points>
<connection>
<GID>86</GID>
<name>N_in2</name></connection>
<intersection>-133.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>975,-133.5,1047.5,-133.5</points>
<connection>
<GID>32</GID>
<name>IN_2</name></connection>
<intersection>975 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>865.5,47.5,869.5,47.5</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<connection>
<GID>188</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>908.5,-102.5,908.5,13</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>900.5,13,908.5,13</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>908.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>863.5,35,863.5,45.5</points>
<intersection>35 1</intersection>
<intersection>38.5 2</intersection>
<intersection>45.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>863.5,35,869,35</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>863.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>863.5,38.5,869.5,38.5</points>
<connection>
<GID>190</GID>
<name>IN_2</name></connection>
<intersection>863.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>863.5,45.5,869.5,45.5</points>
<connection>
<GID>188</GID>
<name>IN_2</name></connection>
<intersection>863.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>886,49,894.5,49</points>
<connection>
<GID>184</GID>
<name>OUT</name></connection>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>888.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>888.5,43.5,888.5,49</points>
<intersection>43.5 4</intersection>
<intersection>49 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>877,43.5,888.5,43.5</points>
<intersection>877 5</intersection>
<intersection>888.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>877,41,877,43.5</points>
<intersection>41 9</intersection>
<intersection>43.5 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>877,41,880,41</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>877 5</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>910.5,-102.5,910.5,49</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>900.5,49,910.5,49</points>
<connection>
<GID>196</GID>
<name>OUT</name></connection>
<intersection>910.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>813,-73.5,820.5,-73.5</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>813 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>813,-75.5,813,-73.5</points>
<connection>
<GID>202</GID>
<name>OUT</name></connection>
<intersection>-73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>813,-83.5,820.5,-83.5</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>813 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>813,-83.5,813,-82.5</points>
<connection>
<GID>204</GID>
<name>OUT</name></connection>
<intersection>-83.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>804.5,-80.5,804.5,-64.5</points>
<intersection>-80.5 1</intersection>
<intersection>-73.5 12</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>804.5,-80.5,807,-80.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>804.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>778.5,-64.5,1031,-64.5</points>
<intersection>778.5 61</intersection>
<intersection>804.5 0</intersection>
<intersection>827 5</intersection>
<intersection>869 17</intersection>
<intersection>890.5 22</intersection>
<intersection>931 31</intersection>
<intersection>957.5 36</intersection>
<intersection>999 45</intersection>
<intersection>1031 60</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>827,-72.5,827,-64.5</points>
<intersection>-72.5 7</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>827,-72.5,895.5,-72.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>827 5</intersection>
<intersection>890.5 22</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>804.5,-73.5,807,-73.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>804.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>869,-82,869,-64.5</points>
<intersection>-82 18</intersection>
<intersection>-75 29</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>869,-82,871.5,-82</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>869 17</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>890.5,-72.5,890.5,-64.5</points>
<intersection>-72.5 7</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>869,-75,871.5,-75</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>869 17</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>931,-78,931,-64.5</points>
<intersection>-78 32</intersection>
<intersection>-71 43</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>931,-78,936,-78</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>931 31</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>957.5,-68.5,957.5,-64.5</points>
<intersection>-68.5 38</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>38</ID>
<points>957.5,-68.5,962.5,-68.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>957.5 36</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>931,-71,936,-71</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>931 31</intersection></hsegment>
<vsegment>
<ID>45</ID>
<points>999,-76.5,999,-64.5</points>
<intersection>-76.5 46</intersection>
<intersection>-69.5 57</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>999,-76.5,1001.5,-76.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>999 45</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>999,-69.5,1001.5,-69.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>999 45</intersection></hsegment>
<vsegment>
<ID>60</ID>
<points>1031,-68,1031,-64.5</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>-64.5 2</intersection></vsegment>
<vsegment>
<ID>61</ID>
<points>778.5,-91.5,778.5,-64.5</points>
<connection>
<GID>28</GID>
<name>OUT_3</name></connection>
<intersection>-64.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>972,-102,972,-70.5</points>
<connection>
<GID>63</GID>
<name>IN_3</name></connection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>968.5,-70.5,972,-70.5</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<intersection>972 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>804,-75.5,807,-75.5</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<connection>
<GID>202</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>793.5,-96,1023.5,-96</points>
<intersection>793.5 5</intersection>
<intersection>814 6</intersection>
<intersection>830.5 3</intersection>
<intersection>892.5 8</intersection>
<intersection>960 17</intersection>
<intersection>1023.5 24</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>830.5,-96,830.5,-76.5</points>
<intersection>-96 1</intersection>
<intersection>-76.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>830.5,-76.5,833.5,-76.5</points>
<connection>
<GID>210</GID>
<name>IN_2</name></connection>
<intersection>830.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>793.5,-151.5,793.5,29.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>-96 1</intersection>
<intersection>-52 29</intersection>
<intersection>-8.5 56</intersection>
<intersection>29.5 77</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>814,-96,814,-88</points>
<intersection>-96 1</intersection>
<intersection>-88 120</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>892.5,-96,892.5,-76.5</points>
<intersection>-96 1</intersection>
<intersection>-89.5 9</intersection>
<intersection>-76.5 12</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>877,-89.5,892.5,-89.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>892.5 8</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>892.5,-76.5,895.5,-76.5</points>
<connection>
<GID>224</GID>
<name>IN_2</name></connection>
<intersection>892.5 8</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>960,-96,960,-72.5</points>
<intersection>-96 1</intersection>
<intersection>-84.5 123</intersection>
<intersection>-72.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>960,-72.5,962.5,-72.5</points>
<connection>
<GID>265</GID>
<name>IN_2</name></connection>
<intersection>960 17</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>1023.5,-96,1023.5,-72</points>
<intersection>-96 1</intersection>
<intersection>-84.5 123</intersection>
<intersection>-72 25</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>1023.5,-72,1031,-72</points>
<connection>
<GID>311</GID>
<name>IN_2</name></connection>
<intersection>1023.5 24</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>793.5,-52,1024.5,-52</points>
<intersection>793.5 5</intersection>
<intersection>816.5 34</intersection>
<intersection>830.5 31</intersection>
<intersection>891 36</intersection>
<intersection>959.5 45</intersection>
<intersection>1024.5 49</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>830.5,-52,830.5,-32.5</points>
<intersection>-52 29</intersection>
<intersection>-32.5 32</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>830.5,-32.5,833,-32.5</points>
<connection>
<GID>106</GID>
<name>IN_2</name></connection>
<intersection>830.5 31</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>816.5,-52,816.5,-46</points>
<intersection>-52 29</intersection>
<intersection>-46 119</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>891,-52,891,-30.5</points>
<intersection>-52 29</intersection>
<intersection>-44 37</intersection>
<intersection>-30.5 40</intersection></vsegment>
<hsegment>
<ID>37</ID>
<points>876,-44,891,-44</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>891 36</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>891,-30.5,895,-30.5</points>
<connection>
<GID>162</GID>
<name>IN_2</name></connection>
<intersection>891 36</intersection></hsegment>
<vsegment>
<ID>45</ID>
<points>959.5,-52,959.5,-28</points>
<intersection>-52 29</intersection>
<intersection>-42 122</intersection>
<intersection>-28 46</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>959.5,-28,961.5,-28</points>
<connection>
<GID>253</GID>
<name>IN_2</name></connection>
<intersection>959.5 45</intersection></hsegment>
<vsegment>
<ID>49</ID>
<points>1024.5,-52,1024.5,-30.5</points>
<intersection>-52 29</intersection>
<intersection>-44.5 50</intersection>
<intersection>-30.5 53</intersection></vsegment>
<hsegment>
<ID>50</ID>
<points>1006.5,-44.5,1024.5,-44.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>1024.5 49</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>1024.5,-30.5,1030.5,-30.5</points>
<connection>
<GID>303</GID>
<name>IN_2</name></connection>
<intersection>1024.5 49</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>793.5,-8.5,1028,-8.5</points>
<intersection>793.5 5</intersection>
<intersection>813.5 61</intersection>
<intersection>830.5 58</intersection>
<intersection>891 63</intersection>
<intersection>945 74</intersection>
<intersection>959 72</intersection>
<intersection>1028 96</intersection></hsegment>
<vsegment>
<ID>58</ID>
<points>830.5,-8.5,830.5,10.5</points>
<intersection>-8.5 56</intersection>
<intersection>10.5 59</intersection></vsegment>
<hsegment>
<ID>59</ID>
<points>830.5,10.5,832.5,10.5</points>
<connection>
<GID>59</GID>
<name>IN_2</name></connection>
<intersection>830.5 58</intersection></hsegment>
<vsegment>
<ID>61</ID>
<points>813.5,-8.5,813.5,-2</points>
<intersection>-8.5 56</intersection>
<intersection>-2 118</intersection></vsegment>
<vsegment>
<ID>63</ID>
<points>891,-8.5,891,11</points>
<intersection>-8.5 56</intersection>
<intersection>-2 64</intersection>
<intersection>11 67</intersection></vsegment>
<hsegment>
<ID>64</ID>
<points>875.5,-2,891,-2</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>891 63</intersection></hsegment>
<hsegment>
<ID>67</ID>
<points>891,11,894.5,11</points>
<connection>
<GID>145</GID>
<name>IN_2</name></connection>
<intersection>891 63</intersection></hsegment>
<vsegment>
<ID>72</ID>
<points>959,-8.5,959,9</points>
<intersection>-8.5 56</intersection>
<intersection>9 73</intersection></vsegment>
<hsegment>
<ID>73</ID>
<points>959,9,961,9</points>
<connection>
<GID>243</GID>
<name>IN_2</name></connection>
<intersection>959 72</intersection></hsegment>
<vsegment>
<ID>74</ID>
<points>945,-8.5,945,-4</points>
<intersection>-8.5 56</intersection>
<intersection>-4 121</intersection></vsegment>
<hsegment>
<ID>77</ID>
<points>793.5,29.5,1028,29.5</points>
<intersection>793.5 5</intersection>
<intersection>811 82</intersection>
<intersection>829.5 79</intersection>
<intersection>890 84</intersection>
<intersection>957.5 90</intersection>
<intersection>1028 105</intersection></hsegment>
<vsegment>
<ID>79</ID>
<points>829.5,29.5,829.5,49.5</points>
<intersection>29.5 77</intersection>
<intersection>49.5 80</intersection></vsegment>
<hsegment>
<ID>80</ID>
<points>829.5,49.5,832,49.5</points>
<connection>
<GID>178</GID>
<name>IN_2</name></connection>
<intersection>829.5 79</intersection></hsegment>
<vsegment>
<ID>82</ID>
<points>811,29.5,811,37</points>
<intersection>29.5 77</intersection>
<intersection>37 117</intersection></vsegment>
<vsegment>
<ID>84</ID>
<points>890,29.5,890,47</points>
<intersection>29.5 77</intersection>
<intersection>35 85</intersection>
<intersection>47 88</intersection></vsegment>
<hsegment>
<ID>85</ID>
<points>875,35,890,35</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>890 84</intersection></hsegment>
<hsegment>
<ID>88</ID>
<points>890,47,894.5,47</points>
<connection>
<GID>196</GID>
<name>IN_2</name></connection>
<intersection>890 84</intersection></hsegment>
<vsegment>
<ID>90</ID>
<points>957.5,29.5,957.5,48</points>
<intersection>29.5 77</intersection>
<intersection>37 91</intersection>
<intersection>48 94</intersection></vsegment>
<hsegment>
<ID>91</ID>
<points>939.5,37,1028,37</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>939.5 125</intersection>
<intersection>957.5 90</intersection>
<intersection>1028 105</intersection></hsegment>
<hsegment>
<ID>94</ID>
<points>957.5,48,961.5,48</points>
<connection>
<GID>232</GID>
<name>IN_2</name></connection>
<intersection>957.5 90</intersection></hsegment>
<vsegment>
<ID>96</ID>
<points>1028,-8.5,1028,8</points>
<intersection>-8.5 56</intersection>
<intersection>-4 97</intersection>
<intersection>8 100</intersection></vsegment>
<hsegment>
<ID>97</ID>
<points>1007,-4,1028,-4</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>1028 96</intersection></hsegment>
<hsegment>
<ID>100</ID>
<points>1028,8,1031.5,8</points>
<connection>
<GID>287</GID>
<name>IN_2</name></connection>
<intersection>1028 96</intersection></hsegment>
<vsegment>
<ID>105</ID>
<points>1028,29.5,1028,52</points>
<intersection>29.5 77</intersection>
<intersection>37 91</intersection>
<intersection>52 106</intersection></vsegment>
<hsegment>
<ID>106</ID>
<points>1028,52,1031.5,52</points>
<connection>
<GID>274</GID>
<name>IN_2</name></connection>
<intersection>1028 105</intersection></hsegment>
<hsegment>
<ID>117</ID>
<points>809.5,37,811,37</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>811 82</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>812.5,-2,813.5,-2</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>813.5 61</intersection></hsegment>
<hsegment>
<ID>119</ID>
<points>815.5,-46,816.5,-46</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>816.5 34</intersection></hsegment>
<hsegment>
<ID>120</ID>
<points>813,-88,814,-88</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>814 6</intersection></hsegment>
<hsegment>
<ID>121</ID>
<points>942,-4,945,-4</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>945 74</intersection></hsegment>
<hsegment>
<ID>122</ID>
<points>942,-42,959.5,-42</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>959.5 45</intersection></hsegment>
<hsegment>
<ID>123</ID>
<points>941.5,-84.5,1023.5,-84.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>941.5 127</intersection>
<intersection>960 17</intersection>
<intersection>1023.5 24</intersection></hsegment>
<vsegment>
<ID>125</ID>
<points>939.5,36,939.5,37</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>37 91</intersection></vsegment>
<vsegment>
<ID>127</ID>
<points>941.5,-85.5,941.5,-84.5</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>-84.5 123</intersection></vsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>803,-88,803,-77.5</points>
<intersection>-88 1</intersection>
<intersection>-84.5 2</intersection>
<intersection>-77.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>803,-88,807,-88</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<intersection>803 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>803,-84.5,807,-84.5</points>
<connection>
<GID>204</GID>
<name>IN_2</name></connection>
<intersection>803 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>803,-77.5,807,-77.5</points>
<connection>
<GID>202</GID>
<name>IN_2</name></connection>
<intersection>803 0</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>826.5,-74.5,833.5,-74.5</points>
<connection>
<GID>199</GID>
<name>OUT</name></connection>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<intersection>828 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>828,-79.5,828,-74.5</points>
<intersection>-79.5 4</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>816,-79.5,828,-79.5</points>
<intersection>816 5</intersection>
<intersection>828 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>816,-81.5,816,-79.5</points>
<intersection>-81.5 9</intersection>
<intersection>-79.5 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>816,-81.5,820.5,-81.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>816 5</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>974,-102,974,-26</points>
<connection>
<GID>63</GID>
<name>IN_2</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>967.5,-26,974,-26</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<intersection>974 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>877.5,-74.5,882.5,-74.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>877.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>877.5,-77,877.5,-74.5</points>
<connection>
<GID>216</GID>
<name>OUT</name></connection>
<intersection>-74.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>877.5,-85.5,882.5,-85.5</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>877.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>877.5,-85.5,877.5,-84</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<intersection>-85.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>976,-102,976,11</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>967,11,976,11</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<intersection>976 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>978,-102,978,50</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>967.5,50,978,50</points>
<connection>
<GID>232</GID>
<name>OUT</name></connection>
<intersection>978 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>865.5,-77,871.5,-77</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<connection>
<GID>216</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1040.5,-102,1040.5,-70</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1037,-70,1040.5,-70</points>
<connection>
<GID>311</GID>
<name>OUT</name></connection>
<intersection>1040.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>864,-89.5,864,-79</points>
<intersection>-89.5 1</intersection>
<intersection>-86 2</intersection>
<intersection>-79 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>864,-89.5,871,-89.5</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<intersection>864 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>864,-86,871.5,-86</points>
<connection>
<GID>218</GID>
<name>IN_2</name></connection>
<intersection>864 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>864,-79,871.5,-79</points>
<connection>
<GID>216</GID>
<name>IN_2</name></connection>
<intersection>864 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>888.5,-74.5,895.5,-74.5</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>888.5 16</intersection>
<intersection>890.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>890.5,-80.5,890.5,-74.5</points>
<intersection>-80.5 4</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>879.5,-80.5,890.5,-80.5</points>
<intersection>879.5 5</intersection>
<intersection>890.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>879.5,-83.5,879.5,-80.5</points>
<intersection>-83.5 9</intersection>
<intersection>-80.5 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>879.5,-83.5,882.5,-83.5</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>879.5 5</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>888.5,-75.5,888.5,-74.5</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>-74.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>888.5,-84.5,889.5,-84.5</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>889.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>889.5,-84.5,889.5,-79</points>
<intersection>-84.5 1</intersection>
<intersection>-79 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>879.5,-79,889.5,-79</points>
<intersection>879.5 5</intersection>
<intersection>889.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>879.5,-79,879.5,-76.5</points>
<intersection>-79 4</intersection>
<intersection>-76.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>879.5,-76.5,882.5,-76.5</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>879.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1042.5,-102,1042.5,-28.5</points>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1036.5,-28.5,1042.5,-28.5</points>
<connection>
<GID>303</GID>
<name>OUT</name></connection>
<intersection>1042.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>940.5,51,946.5,51</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>940.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>940.5,48.5,940.5,51</points>
<connection>
<GID>228</GID>
<name>OUT</name></connection>
<intersection>51 1</intersection></vsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>940.5,40,946.5,40</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<intersection>940.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>940.5,40,940.5,41.5</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<intersection>40 1</intersection></vsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1044.5,-102,1044.5,10</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1037.5,10,1044.5,10</points>
<connection>
<GID>287</GID>
<name>OUT</name></connection>
<intersection>1044.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>741,-97.5,741,-58.5</points>
<intersection>-97.5 1</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>738,-97.5,741,-97.5</points>
<connection>
<GID>288</GID>
<name>OUT</name></connection>
<intersection>741 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>738.5,-58.5,744.5,-58.5</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>738.5 3</intersection>
<intersection>741 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>738.5,-58.5,738.5,21.5</points>
<intersection>-58.5 2</intersection>
<intersection>21.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>738.5,21.5,798.5,21.5</points>
<intersection>738.5 3</intersection>
<intersection>781.5 6</intersection>
<intersection>798.5 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>781.5,4,781.5,21.5</points>
<intersection>4 7</intersection>
<intersection>21.5 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>781.5,4,807,4</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>781.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>798.5,11,798.5,21.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>21.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>929.5,48.5,934.5,48.5</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<connection>
<GID>228</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1046.5,-102,1046.5,54</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1037.5,54,1046.5,54</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<intersection>1046.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>927.5,36,927.5,46.5</points>
<intersection>36 1</intersection>
<intersection>39.5 2</intersection>
<intersection>46.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>927.5,36,933.5,36</points>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection>
<intersection>927.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>927.5,39.5,934.5,39.5</points>
<connection>
<GID>229</GID>
<name>IN_2</name></connection>
<intersection>927.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>927.5,46.5,934.5,46.5</points>
<connection>
<GID>228</GID>
<name>IN_2</name></connection>
<intersection>927.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>952.5,50,961.5,50</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<connection>
<GID>226</GID>
<name>OUT</name></connection>
<intersection>953.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>953.5,44,953.5,50</points>
<intersection>44 4</intersection>
<intersection>50 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>942.5,44,953.5,44</points>
<intersection>942.5 5</intersection>
<intersection>953.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>942.5,42,942.5,44</points>
<intersection>42 9</intersection>
<intersection>44 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>942.5,42,946.5,42</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>942.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>952.5,41,954.5,41</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<intersection>954.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>954.5,41,954.5,46</points>
<intersection>41 1</intersection>
<intersection>46 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>942.5,46,954.5,46</points>
<intersection>942.5 5</intersection>
<intersection>954.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>942.5,46,942.5,49</points>
<intersection>46 4</intersection>
<intersection>49 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>942.5,49,946.5,49</points>
<connection>
<GID>226</GID>
<name>IN_1</name></connection>
<intersection>942.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1043.5,-132.5,1043.5,-109</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<connection>
<GID>98</GID>
<name>N_in3</name></connection>
<intersection>-132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1043.5,-132.5,1047.5,-132.5</points>
<connection>
<GID>32</GID>
<name>IN_3</name></connection>
<intersection>1043.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>942.5,12,948.5,12</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>942.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>942.5,8.5,942.5,12</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<intersection>12 1</intersection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>942.5,0.5,948.5,0.5</points>
<connection>
<GID>235</GID>
<name>IN_1</name></connection>
<intersection>942.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>942.5,0.5,942.5,1.5</points>
<connection>
<GID>237</GID>
<name>OUT</name></connection>
<intersection>0.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>907.5,-115,907.5,-109.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<connection>
<GID>76</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>929.5,8.5,936.5,8.5</points>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection>
<connection>
<GID>236</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>846,-115,846,-109</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<connection>
<GID>70</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>927,-4,927,6.5</points>
<intersection>-4 1</intersection>
<intersection>-0.5 2</intersection>
<intersection>6.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>927,-4,936,-4</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<intersection>927 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>927,-0.5,936.5,-0.5</points>
<connection>
<GID>237</GID>
<name>IN_2</name></connection>
<intersection>927 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>927,6.5,936.5,6.5</points>
<connection>
<GID>236</GID>
<name>IN_2</name></connection>
<intersection>927 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>954.5,11,961,11</points>
<connection>
<GID>234</GID>
<name>OUT</name></connection>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>957.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>957.5,5,957.5,11</points>
<intersection>5 4</intersection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>944.5,5,957.5,5</points>
<intersection>944.5 5</intersection>
<intersection>957.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>944.5,2.5,944.5,5</points>
<intersection>2.5 6</intersection>
<intersection>5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>944.5,2.5,948.5,2.5</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>944.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>954.5,1.5,955.5,1.5</points>
<connection>
<GID>235</GID>
<name>OUT</name></connection>
<intersection>955.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>955.5,1.5,955.5,8</points>
<intersection>1.5 1</intersection>
<intersection>8 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>944.5,8,955.5,8</points>
<intersection>944.5 5</intersection>
<intersection>955.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>944.5,8,944.5,10</points>
<intersection>8 4</intersection>
<intersection>10 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>944.5,10,948.5,10</points>
<connection>
<GID>234</GID>
<name>IN_1</name></connection>
<intersection>944.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>975,-115,975,-109</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<connection>
<GID>86</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>942.5,-25.5,948,-25.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>942.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>942.5,-29.5,942.5,-25.5</points>
<connection>
<GID>249</GID>
<name>OUT</name></connection>
<intersection>-25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>942.5,-38,948,-38</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<intersection>942.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>942.5,-38,942.5,-36.5</points>
<connection>
<GID>250</GID>
<name>OUT</name></connection>
<intersection>-38 1</intersection></vsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>927.5,-29.5,936.5,-29.5</points>
<connection>
<GID>251</GID>
<name>OUT_0</name></connection>
<connection>
<GID>249</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>925.5,-42,925.5,-31.5</points>
<intersection>-42 1</intersection>
<intersection>-38.5 2</intersection>
<intersection>-31.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>925.5,-42,936,-42</points>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>925.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>925.5,-38.5,936.5,-38.5</points>
<connection>
<GID>250</GID>
<name>IN_2</name></connection>
<intersection>925.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>925.5,-31.5,936.5,-31.5</points>
<connection>
<GID>249</GID>
<name>IN_2</name></connection>
<intersection>925.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>954,-26,961.5,-26</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<intersection>954 10</intersection>
<intersection>958 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>958,-33.5,958,-26</points>
<intersection>-33.5 4</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>943.5,-33.5,958,-33.5</points>
<intersection>943.5 5</intersection>
<intersection>958 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>943.5,-36,943.5,-33.5</points>
<intersection>-36 6</intersection>
<intersection>-33.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>943.5,-36,948,-36</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>943.5 5</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>954,-26.5,954,-26</points>
<connection>
<GID>247</GID>
<name>OUT</name></connection>
<intersection>-26 1</intersection></vsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>954,-37,957,-37</points>
<connection>
<GID>248</GID>
<name>OUT</name></connection>
<intersection>957 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>957,-37,957,-31</points>
<intersection>-37 1</intersection>
<intersection>-31 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>943.5,-31,957,-31</points>
<intersection>943.5 5</intersection>
<intersection>957 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>943.5,-31,943.5,-27.5</points>
<intersection>-31 4</intersection>
<intersection>-27.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>943.5,-27.5,948,-27.5</points>
<connection>
<GID>247</GID>
<name>IN_1</name></connection>
<intersection>943.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>942,-69.5,947,-69.5</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>942 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>942,-73,942,-69.5</points>
<connection>
<GID>258</GID>
<name>OUT</name></connection>
<intersection>-69.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>942,-81,947,-81</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>942 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>942,-81,942,-80</points>
<connection>
<GID>259</GID>
<name>OUT</name></connection>
<intersection>-81 1</intersection></vsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>926.5,-73,936,-73</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<connection>
<GID>258</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>925.5,-85.5,925.5,-75</points>
<intersection>-85.5 1</intersection>
<intersection>-82 2</intersection>
<intersection>-75 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>925.5,-85.5,935.5,-85.5</points>
<connection>
<GID>263</GID>
<name>OUT_0</name></connection>
<intersection>925.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>925.5,-82,936,-82</points>
<connection>
<GID>259</GID>
<name>IN_2</name></connection>
<intersection>925.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>925.5,-75,936,-75</points>
<connection>
<GID>258</GID>
<name>IN_2</name></connection>
<intersection>925.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>953,-70.5,962.5,-70.5</points>
<connection>
<GID>255</GID>
<name>OUT</name></connection>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<intersection>958.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>958.5,-76,958.5,-70.5</points>
<intersection>-76 4</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>943.5,-76,958.5,-76</points>
<intersection>943.5 5</intersection>
<intersection>958.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>943.5,-79,943.5,-76</points>
<intersection>-79 9</intersection>
<intersection>-76 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>943.5,-79,947,-79</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>943.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>953,-80,956.5,-80</points>
<connection>
<GID>257</GID>
<name>OUT</name></connection>
<intersection>956.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>956.5,-80,956.5,-74</points>
<intersection>-80 1</intersection>
<intersection>-74 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>943.5,-74,956.5,-74</points>
<intersection>943.5 5</intersection>
<intersection>956.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>943.5,-74,943.5,-71.5</points>
<intersection>-74 4</intersection>
<intersection>-71.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>943.5,-71.5,947,-71.5</points>
<connection>
<GID>255</GID>
<name>IN_1</name></connection>
<intersection>943.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1009.5,54.5,1014.5,54.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>1009.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1009.5,50,1009.5,54.5</points>
<connection>
<GID>270</GID>
<name>OUT</name></connection>
<intersection>54.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1009.5,41.5,1014.5,41.5</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<intersection>1009.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>1009.5,41.5,1009.5,42.5</points>
<connection>
<GID>271</GID>
<name>OUT</name></connection>
<intersection>41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>743.5,-91,743.5,-65</points>
<intersection>-91 2</intersection>
<intersection>-65 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>738,-91,743.5,-91</points>
<connection>
<GID>286</GID>
<name>OUT</name></connection>
<intersection>743.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>737.5,-65,744.5,-65</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>737.5 4</intersection>
<intersection>743.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>737.5,-65,737.5,26</points>
<intersection>-65 3</intersection>
<intersection>10.5 6</intersection>
<intersection>26 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>737.5,26,869.5,26</points>
<intersection>737.5 4</intersection>
<intersection>869.5 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>737.5,10.5,858.5,10.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>737.5 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>869.5,3.5,869.5,26</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>26 5</intersection></vsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>995.5,50,1003.5,50</points>
<connection>
<GID>272</GID>
<name>OUT_0</name></connection>
<connection>
<GID>270</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>996,37,996,48</points>
<intersection>37 1</intersection>
<intersection>40.5 2</intersection>
<intersection>48 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>996,37,1003,37</points>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection>
<intersection>996 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>996,40.5,1003.5,40.5</points>
<connection>
<GID>271</GID>
<name>IN_2</name></connection>
<intersection>996 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>996,48,1003.5,48</points>
<connection>
<GID>270</GID>
<name>IN_2</name></connection>
<intersection>996 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1020.5,54,1031.5,54</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>1020.5 13</intersection>
<intersection>1023 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1023,47,1023,54</points>
<intersection>47 4</intersection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1011,47,1023,47</points>
<intersection>1011 5</intersection>
<intersection>1023 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>1011,43.5,1011,47</points>
<intersection>43.5 9</intersection>
<intersection>47 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>1011,43.5,1014.5,43.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>1011 5</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>1020.5,53.5,1020.5,54</points>
<connection>
<GID>268</GID>
<name>OUT</name></connection>
<intersection>54 1</intersection></vsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1020.5,42.5,1025,42.5</points>
<connection>
<GID>269</GID>
<name>OUT</name></connection>
<intersection>1025 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1025,42.5,1025,49</points>
<intersection>42.5 1</intersection>
<intersection>49 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1011,49,1025,49</points>
<intersection>1011 5</intersection>
<intersection>1025 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>1011,49,1011,52.5</points>
<intersection>49 4</intersection>
<intersection>52.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>1011,52.5,1014.5,52.5</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>1011 5</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1007.5,11,1013.5,11</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>1007.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1007.5,8.5,1007.5,11</points>
<connection>
<GID>281</GID>
<name>OUT</name></connection>
<intersection>11 1</intersection></vsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1007.5,1,1013.5,1</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>1007.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>1007.5,1,1007.5,1.5</points>
<connection>
<GID>283</GID>
<name>OUT</name></connection>
<intersection>1 1</intersection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>996,8.5,1001.5,8.5</points>
<connection>
<GID>284</GID>
<name>OUT_0</name></connection>
<connection>
<GID>281</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>994.5,-4,994.5,6.5</points>
<intersection>-4 1</intersection>
<intersection>-0.5 2</intersection>
<intersection>6.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>994.5,-4,1001,-4</points>
<connection>
<GID>285</GID>
<name>OUT_0</name></connection>
<intersection>994.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>994.5,-0.5,1001.5,-0.5</points>
<connection>
<GID>283</GID>
<name>IN_2</name></connection>
<intersection>994.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>994.5,6.5,1001.5,6.5</points>
<connection>
<GID>281</GID>
<name>IN_2</name></connection>
<intersection>994.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1019.5,10,1031.5,10</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<connection>
<GID>287</GID>
<name>IN_1</name></connection>
<intersection>1021.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1021.5,5.5,1021.5,10</points>
<intersection>5.5 4</intersection>
<intersection>10 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1009.5,5.5,1021.5,5.5</points>
<intersection>1009.5 5</intersection>
<intersection>1021.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>1009.5,3,1009.5,5.5</points>
<intersection>3 9</intersection>
<intersection>5.5 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>1009.5,3,1013.5,3</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>1009.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1019.5,2,1020.5,2</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<intersection>1020.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1020.5,2,1020.5,6</points>
<intersection>2 1</intersection>
<intersection>6 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1009.5,6,1020.5,6</points>
<intersection>1009.5 5</intersection>
<intersection>1020.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>1009.5,6,1009.5,9</points>
<intersection>6 4</intersection>
<intersection>9 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>1009.5,9,1013.5,9</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>1009.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1007,-28,1012,-28</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>1007 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1007,-31.5,1007,-28</points>
<connection>
<GID>295</GID>
<name>OUT</name></connection>
<intersection>-28 1</intersection></vsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1007,-41,1012,-41</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<intersection>1007 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>1007,-41,1007,-38.5</points>
<connection>
<GID>297</GID>
<name>OUT</name></connection>
<intersection>-41 1</intersection></vsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>995,-31.5,1001,-31.5</points>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection>
<connection>
<GID>295</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>993,-44.5,993,-33.5</points>
<intersection>-44.5 1</intersection>
<intersection>-40.5 2</intersection>
<intersection>-33.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>993,-44.5,1000.5,-44.5</points>
<connection>
<GID>301</GID>
<name>OUT_0</name></connection>
<intersection>993 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>993,-40.5,1001,-40.5</points>
<connection>
<GID>297</GID>
<name>IN_2</name></connection>
<intersection>993 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>993,-33.5,1001,-33.5</points>
<connection>
<GID>295</GID>
<name>IN_2</name></connection>
<intersection>993 0</intersection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1018,-28.5,1030.5,-28.5</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<intersection>1018 13</intersection>
<intersection>1020 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1020,-35.5,1020,-28.5</points>
<intersection>-35.5 4</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1009,-35.5,1020,-35.5</points>
<intersection>1009 5</intersection>
<intersection>1020 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>1009,-39,1009,-35.5</points>
<intersection>-39 9</intersection>
<intersection>-35.5 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>1009,-39,1012,-39</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>1009 5</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>1018,-29,1018,-28.5</points>
<connection>
<GID>291</GID>
<name>OUT</name></connection>
<intersection>-28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1018,-40,1019,-40</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<intersection>1019 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1019,-40,1019,-34</points>
<intersection>-40 1</intersection>
<intersection>-34 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1009,-34,1019,-34</points>
<intersection>1009 5</intersection>
<intersection>1019 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>1009,-34,1009,-30</points>
<intersection>-34 4</intersection>
<intersection>-30 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>1009,-30,1012,-30</points>
<connection>
<GID>291</GID>
<name>IN_1</name></connection>
<intersection>1009 5</intersection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1007.5,-69,1012,-69</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>1007.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1007.5,-71.5,1007.5,-69</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<intersection>-69 1</intersection></vsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1007.5,-80.5,1012,-80.5</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<intersection>1007.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>1007.5,-80.5,1007.5,-78.5</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<intersection>-80.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>995.5,-71.5,1001.5,-71.5</points>
<connection>
<GID>309</GID>
<name>OUT_0</name></connection>
<connection>
<GID>307</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>994.5,-84.5,994.5,-73.5</points>
<intersection>-84.5 1</intersection>
<intersection>-80.5 2</intersection>
<intersection>-73.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>994.5,-84.5,1001,-84.5</points>
<connection>
<GID>310</GID>
<name>OUT_0</name></connection>
<intersection>994.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>994.5,-80.5,1001.5,-80.5</points>
<connection>
<GID>308</GID>
<name>IN_2</name></connection>
<intersection>994.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>994.5,-73.5,1001.5,-73.5</points>
<connection>
<GID>307</GID>
<name>IN_2</name></connection>
<intersection>994.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1018,-70,1031,-70</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<intersection>1019 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1019,-76,1019,-70</points>
<intersection>-76 4</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1009,-76,1019,-76</points>
<intersection>1009 5</intersection>
<intersection>1019 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>1009,-78.5,1009,-76</points>
<intersection>-78.5 9</intersection>
<intersection>-76 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>1009,-78.5,1012,-78.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>1009 5</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1018,-79.5,1020.5,-79.5</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>1020.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1020.5,-79.5,1020.5,-73.5</points>
<intersection>-79.5 1</intersection>
<intersection>-73.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1009,-73.5,1020.5,-73.5</points>
<intersection>1009 5</intersection>
<intersection>1020.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>1009,-73.5,1009,-71</points>
<intersection>-73.5 4</intersection>
<intersection>-71 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>1009,-71,1012,-71</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>1009 5</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>783.5,-93.5,783.5,18.5</points>
<intersection>-93.5 2</intersection>
<intersection>18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>783.5,18.5,1031.5,18.5</points>
<intersection>783.5 0</intersection>
<intersection>805.5 3</intersection>
<intersection>832.5 5</intersection>
<intersection>866 10</intersection>
<intersection>894.5 12</intersection>
<intersection>934 17</intersection>
<intersection>961 19</intersection>
<intersection>997 21</intersection>
<intersection>1031.5 23</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>778.5,-93.5,783.5,-93.5</points>
<connection>
<GID>28</GID>
<name>OUT_1</name></connection>
<intersection>783.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>805.5,6,805.5,18.5</points>
<intersection>6 7</intersection>
<intersection>13 8</intersection>
<intersection>18.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>832.5,14.5,832.5,18.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>18.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>805.5,6,807,6</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>805.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>805.5,13,807,13</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>805.5 3</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>866,5.5,866,18.5</points>
<intersection>5.5 14</intersection>
<intersection>12.5 15</intersection>
<intersection>18.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>894.5,15,894.5,18.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>18.5 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>866,5.5,869.5,5.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>866 10</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>866,12.5,869.5,12.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>866 10</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>934,3.5,934,18.5</points>
<intersection>3.5 25</intersection>
<intersection>10.5 26</intersection>
<intersection>18.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>961,13,961,18.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>18.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>997,3.5,997,18.5</points>
<intersection>3.5 28</intersection>
<intersection>10.5 29</intersection>
<intersection>18.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>1031.5,12,1031.5,18.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>18.5 1</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>934,3.5,936.5,3.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>934 17</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>934,10.5,936.5,10.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>934 17</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>997,3.5,1001.5,3.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>997 21</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>997,10.5,1001.5,10.5</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>997 21</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>863,-2,863,8.5</points>
<intersection>-2 2</intersection>
<intersection>1.5 4</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>863,8.5,869.5,8.5</points>
<connection>
<GID>128</GID>
<name>IN_2</name></connection>
<intersection>863 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>863,-2,869.5,-2</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>863 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>863,1.5,869.5,1.5</points>
<connection>
<GID>132</GID>
<name>IN_2</name></connection>
<intersection>863 0</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>986.5,-3.5,986.5,1.5</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>986.5,1.5,1001.5,1.5</points>
<connection>
<GID>283</GID>
<name>IN_1</name></connection>
<intersection>986.5 0</intersection>
<intersection>990 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>990,1.5,990,8.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>1.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>919,-3.5,919,1.5</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>919,1.5,936.5,1.5</points>
<connection>
<GID>237</GID>
<name>IN_1</name></connection>
<intersection>919 0</intersection>
<intersection>923.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>923.5,1.5,923.5,8.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>1.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>750.5,-151.5,750.5,-93.5</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>750.5,-93.5,772.5,-93.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>750.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>756.5,-151.5,756.5,-94.5</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<intersection>-94.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>756.5,-94.5,772.5,-94.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>756.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>829.5,-82.5,829.5,-78</points>
<intersection>-82.5 2</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>820.5,-78,829.5,-78</points>
<intersection>820.5 3</intersection>
<intersection>829.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>826.5,-82.5,829.5,-82.5</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>829.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>820.5,-78,820.5,-75.5</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>-78 1</intersection></vsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>887,40,887,45</points>
<intersection>40 2</intersection>
<intersection>45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>880,45,887,45</points>
<intersection>880 3</intersection>
<intersection>887 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>886,40,887,40</points>
<connection>
<GID>186</GID>
<name>OUT</name></connection>
<intersection>887 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>880,45,880,48</points>
<connection>
<GID>184</GID>
<name>IN_1</name></connection>
<intersection>45 1</intersection></vsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>790.5,-117.5,790.5,-32</points>
<intersection>-117.5 1</intersection>
<intersection>-40 4</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>769.5,-117.5,790.5,-117.5</points>
<connection>
<GID>40</GID>
<name>N_in1</name></connection>
<intersection>790.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>790.5,-32,798.5,-32</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>790.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>790.5,-40,809,-40</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>790.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>853,-128,853,-31.5</points>
<intersection>-128 1</intersection>
<intersection>-38.5 4</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>770,-128,853,-128</points>
<connection>
<GID>48</GID>
<name>N_in1</name></connection>
<intersection>853 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>853,-31.5,859,-31.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>853 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>853,-38.5,869.5,-38.5</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>853 0</intersection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>918,-141.5,918,-29.5</points>
<intersection>-141.5 1</intersection>
<intersection>-36.5 6</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>780,-141.5,918,-141.5</points>
<intersection>780 3</intersection>
<intersection>918 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>918,-29.5,921.5,-29.5</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>918 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>780,-141.5,780,-138.5</points>
<intersection>-141.5 1</intersection>
<intersection>-138.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>770,-138.5,780,-138.5</points>
<connection>
<GID>53</GID>
<name>N_in1</name></connection>
<intersection>780 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>918,-36.5,936.5,-36.5</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<intersection>918 0</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>985,-47.5,985,-31.5</points>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection>
<intersection>-38.5 1</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>985,-38.5,1001,-38.5</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>985 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>985,-31.5,989,-31.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>985 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>841.5,-58.5,841.5,-12.5</points>
<intersection>-58.5 2</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>768.5,-12.5,841.5,-12.5</points>
<intersection>768.5 4</intersection>
<intersection>841.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>841.5,-58.5,920.5,-58.5</points>
<intersection>841.5 0</intersection>
<intersection>920.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>920.5,-80,920.5,-58.5</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>-80 5</intersection>
<intersection>-58.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>768.5,-12.5,768.5,3.5</points>
<connection>
<GID>50</GID>
<name>N_in1</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>920.5,-80,936,-80</points>
<connection>
<GID>259</GID>
<name>IN_1</name></connection>
<intersection>920.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>988,-80.5,988,-78.5</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>988,-78.5,1001.5,-78.5</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>988 0</intersection>
<intersection>989.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>989.5,-78.5,989.5,-71.5</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>-78.5 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>620.561,145.494,1844.56,-459.506</PageViewport>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>648,-49</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>184.5,-45.5</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>648,-57</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>177,-45.5</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_TOGGLE</type>
<position>169.5,-45.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>648,-64</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_TOGGLE</type>
<position>162,-45.5</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_TOGGLE</type>
<position>648,-72</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>161,-42</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>746,-60</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>108 </input>
<input>
<ID>IN_3</ID>107 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>169.5,-41.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>177,-41.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_TOGGLE</type>
<position>659,-30.5</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>184.5,-41.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_TOGGLE</type>
<position>662,-30.5</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_TOGGLE</type>
<position>665,-30.5</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_TOGGLE</type>
<position>668,-30.5</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_AND2</type>
<position>668,-47.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_AND2</type>
<position>667.5,-56</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_AND2</type>
<position>667.5,-63.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND2</type>
<position>668,-71</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>105</ID>
<type>AI_XOR2</type>
<position>681,-47</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>AI_XOR2</type>
<position>681,-54.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AI_XOR2</type>
<position>681,-62.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>AI_XOR2</type>
<position>681,-70</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AI_XOR2</type>
<position>696.5,-46.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AI_XOR2</type>
<position>697,-55</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>AI_XOR2</type>
<position>697,-63</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_AND3</type>
<position>220,-57</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>69 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_INVERTER</type>
<position>205.5,-62</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>134</ID>
<type>AI_XOR2</type>
<position>697,-70.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_INVERTER</type>
<position>199,-64.5</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_AND2</type>
<position>213,-71.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>AI_XOR2</type>
<position>714,-47</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_AND3</type>
<position>213,-78.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>71 </input>
<input>
<ID>IN_2</ID>69 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>141</ID>
<type>AE_OR3</type>
<position>237,-70.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>60 </input>
<input>
<ID>IN_2</ID>61 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>142</ID>
<type>AI_XOR2</type>
<position>714,-55.5</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>AI_XOR2</type>
<position>714,-63.5</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>102 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>AI_XOR2</type>
<position>714,-71</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_OR2</type>
<position>60.5,-57</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND2</type>
<position>231,-88</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_AND3</type>
<position>213,-107.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>74 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_AND2</type>
<position>213,-114</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AE_OR3</type>
<position>233.5,-107</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>65 </input>
<input>
<ID>IN_2</ID>66 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_INVERTER</type>
<position>204,-72.5</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_INVERTER</type>
<position>207,-76.5</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_INVERTER</type>
<position>206.5,-98</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_INVERTER</type>
<position>207,-109.5</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_INVERTER</type>
<position>207,-115</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>252,-70</position>
<input>
<ID>N_in0</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>GA_LED</type>
<position>252,-87.5</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>GA_LED</type>
<position>252.5,-104.5</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AO_XNOR2</type>
<position>202.5,-85.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>71 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AO_XNOR2</type>
<position>202.5,-91.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_AND3</type>
<position>217.5,-98.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>84 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_INVERTER</type>
<position>209,-102</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>657.5,-49,657.5,-48.5</points>
<intersection>-49 2</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>657.5,-48.5,665,-48.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>657.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>650,-49,657.5,-49</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>657.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>662,-70,662,-32.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<intersection>-70 7</intersection>
<intersection>-62.5 5</intersection>
<intersection>-55 3</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>662,-46.5,665,-46.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>662 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>662,-55,664.5,-55</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>662 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>662,-62.5,664.5,-62.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>662 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>662,-70,665,-70</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>662 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>650,-57,664.5,-57</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>657,-64.5,657,-64</points>
<intersection>-64.5 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>650,-64,657,-64</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>657 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>657,-64.5,664.5,-64.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>657 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>650,-72,665,-72</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<connection>
<GID>103</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>659,-43,659,-32.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>659,-43,676.5,-43</points>
<intersection>659 0</intersection>
<intersection>676.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>676.5,-69,676.5,-43</points>
<intersection>-69 9</intersection>
<intersection>-61.5 7</intersection>
<intersection>-53.5 5</intersection>
<intersection>-46 3</intersection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>676.5,-46,678,-46</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>676.5 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>676.5,-53.5,678,-53.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>676.5 2</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>676.5,-61.5,678,-61.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>676.5 2</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>676.5,-69,678,-69</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>676.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>674.5,-48,674.5,-47.5</points>
<intersection>-48 1</intersection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>674.5,-48,678,-48</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>674.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>671,-47.5,674.5,-47.5</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>674.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206,-64.5,206,-57</points>
<intersection>-64.5 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206,-57,217,-57</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>206 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>202,-64.5,206,-64.5</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<intersection>206 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-68.5,225,-57</points>
<intersection>-68.5 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,-68.5,234,-68.5</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,-57,225,-57</points>
<connection>
<GID>131</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-71.5,225,-70.5</points>
<intersection>-71.5 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,-70.5,234,-70.5</points>
<connection>
<GID>141</GID>
<name>IN_1</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-71.5,225,-71.5</points>
<connection>
<GID>137</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-78.5,225,-72.5</points>
<intersection>-78.5 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,-72.5,234,-72.5</points>
<connection>
<GID>141</GID>
<name>IN_2</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-78.5,225,-78.5</points>
<connection>
<GID>139</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>674,-56,674,-55.5</points>
<intersection>-56 1</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>670.5,-56,674,-56</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<intersection>674 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>674,-55.5,678,-55.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>674 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>670.5,-63.5,678,-63.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<connection>
<GID>109</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>671,-71,678,-71</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<connection>
<GID>111</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223,-107.5,223,-107</points>
<intersection>-107.5 2</intersection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223,-107,230.5,-107</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>223 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-107.5,223,-107.5</points>
<connection>
<GID>153</GID>
<name>OUT</name></connection>
<intersection>223 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223,-114,223,-109</points>
<intersection>-114 2</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223,-109,230.5,-109</points>
<connection>
<GID>157</GID>
<name>IN_2</name></connection>
<intersection>223 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-114,223,-114</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<intersection>223 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-62,177,-47.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,-62,202.5,-62</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>177 0</intersection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-72.5,192,-62</points>
<intersection>-72.5 3</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-72.5,201,-72.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>176 4</intersection>
<intersection>180.5 10</intersection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>176,-113,176,-72.5</points>
<intersection>-113 9</intersection>
<intersection>-105.5 7</intersection>
<intersection>-72.5 3</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>176,-105.5,210,-105.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>176 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>176,-113,210,-113</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>176 4</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>180.5,-84.5,180.5,-72.5</points>
<intersection>-84.5 11</intersection>
<intersection>-72.5 3</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>180.5,-84.5,199.5,-84.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>180.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-107.5,162,-47.5</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<intersection>-107.5 9</intersection>
<intersection>-98.5 7</intersection>
<intersection>-76.5 3</intersection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162,-64.5,196,-64.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>162,-76.5,204,-76.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>162,-98.5,164,-98.5</points>
<intersection>162 0</intersection>
<intersection>164 10</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>162,-107.5,210,-107.5</points>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<intersection>162 0</intersection>
<intersection>196 12</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>164,-98.5,164,-90.5</points>
<intersection>-98.5 7</intersection>
<intersection>-90.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>164,-90.5,199.5,-90.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>164 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>196,-107.5,196,-96.5</points>
<intersection>-107.5 9</intersection>
<intersection>-96.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>196,-96.5,214.5,-96.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>196 12</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-109.5,169.5,-47.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 9</intersection>
<intersection>-102.5 7</intersection>
<intersection>-80.5 3</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-59,217,-59</points>
<connection>
<GID>131</GID>
<name>IN_2</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>169.5,-80.5,210,-80.5</points>
<connection>
<GID>139</GID>
<name>IN_2</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>169.5,-102.5,193,-102.5</points>
<intersection>169.5 0</intersection>
<intersection>193 10</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>169.5,-109.5,204,-109.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection>
<intersection>201.5 12</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>193,-102.5,193,-92.5</points>
<intersection>-102.5 7</intersection>
<intersection>-92.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>193,-92.5,199.5,-92.5</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>193 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>201.5,-109.5,201.5,-102</points>
<intersection>-109.5 9</intersection>
<intersection>-102 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>201.5,-102,206,-102</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>201.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>207,-72.5,210,-72.5</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-115,184.5,-47.5</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>-115 9</intersection>
<intersection>-98 7</intersection>
<intersection>-78.5 3</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,-70.5,210,-70.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>184.5,-78.5,210,-78.5</points>
<connection>
<GID>139</GID>
<name>IN_1</name></connection>
<intersection>184.5 0</intersection>
<intersection>186.5 10</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>184.5,-98,203.5,-98</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>184.5,-115,204,-115</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>186.5,-86.5,186.5,-78.5</points>
<intersection>-86.5 11</intersection>
<intersection>-78.5 3</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>186.5,-86.5,199.5,-86.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>186.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-76.5,210,-76.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,-71.5,689,-70</points>
<intersection>-71.5 1</intersection>
<intersection>-70 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>689,-71.5,694,-71.5</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>689 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>684,-70,689,-70</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>689 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-109.5,210,-109.5</points>
<connection>
<GID>153</GID>
<name>IN_2</name></connection>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-115,210,-115</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-70.5,245.5,-70</points>
<intersection>-70.5 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245.5,-70,251,-70</points>
<connection>
<GID>169</GID>
<name>N_in0</name></connection>
<intersection>245.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>240,-70.5,245.5,-70.5</points>
<connection>
<GID>141</GID>
<name>OUT</name></connection>
<intersection>245.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242.5,-88,242.5,-87.5</points>
<intersection>-88 2</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242.5,-87.5,251,-87.5</points>
<connection>
<GID>171</GID>
<name>N_in0</name></connection>
<intersection>242.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234,-88,242.5,-88</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>242.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-107,244,-104.5</points>
<intersection>-107 2</intersection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,-104.5,251.5,-104.5</points>
<connection>
<GID>173</GID>
<name>N_in0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>236.5,-107,244,-107</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216.5,-87,216.5,-85.5</points>
<intersection>-87 1</intersection>
<intersection>-85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216.5,-87,228,-87</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>216.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>205.5,-85.5,216.5,-85.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>216.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216.5,-91.5,216.5,-89</points>
<intersection>-91.5 1</intersection>
<intersection>-89 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205.5,-91.5,216.5,-91.5</points>
<connection>
<GID>177</GID>
<name>OUT</name></connection>
<intersection>216.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216.5,-89,228,-89</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>216.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>208.5,-55,217,-55</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>208.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>208.5,-62,208.5,-55</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>-55 1</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,-105,225.5,-98.5</points>
<intersection>-105 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225.5,-105,230.5,-105</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,-98.5,225.5,-98.5</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,-98.5,212,-98</points>
<intersection>-98.5 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209.5,-98,212,-98</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>212,-98.5,214.5,-98.5</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>212 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-102,213,-100.5</points>
<intersection>-102 2</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213,-100.5,214.5,-100.5</points>
<connection>
<GID>179</GID>
<name>IN_2</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>212,-102,213,-102</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,-64,689,-62.5</points>
<intersection>-64 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>684,-62.5,689,-62.5</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>689 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>689,-64,694,-64</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>689 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,-56,689,-54.5</points>
<intersection>-56 2</intersection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>684,-54.5,689,-54.5</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>689 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>689,-56,694,-56</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>689 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>688.5,-47.5,688.5,-47</points>
<intersection>-47.5 2</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>684,-47,688.5,-47</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<intersection>688.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>688.5,-47.5,693.5,-47.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>688.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>665,-42,665,-32.5</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>665,-42,691.5,-42</points>
<intersection>665 0</intersection>
<intersection>691.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>691.5,-69.5,691.5,-42</points>
<intersection>-69.5 9</intersection>
<intersection>-62 7</intersection>
<intersection>-54 5</intersection>
<intersection>-45.5 3</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>691.5,-45.5,693.5,-45.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>691.5 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>691.5,-54,694,-54</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>691.5 2</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>691.5,-62,694,-62</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>691.5 2</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>691.5,-69.5,694,-69.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>691.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>705,-48,705,-46.5</points>
<intersection>-48 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>705,-48,711,-48</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>705 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>699.5,-46.5,705,-46.5</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>705 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>705.5,-56.5,705.5,-55</points>
<intersection>-56.5 1</intersection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>705.5,-56.5,711,-56.5</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>705.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>700,-55,705.5,-55</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<intersection>705.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>705.5,-64.5,705.5,-63</points>
<intersection>-64.5 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>705.5,-64.5,711,-64.5</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>705.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>700,-63,705.5,-63</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<intersection>705.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>705.5,-72,705.5,-70.5</points>
<intersection>-72 1</intersection>
<intersection>-70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>705.5,-72,711,-72</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>705.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>700,-70.5,705.5,-70.5</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<intersection>705.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668,-41,668,-32.5</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>668,-41,709,-41</points>
<intersection>668 0</intersection>
<intersection>709 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>709,-70,709,-41</points>
<intersection>-70 9</intersection>
<intersection>-62.5 7</intersection>
<intersection>-54.5 5</intersection>
<intersection>-46 3</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>709,-46,711,-46</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>709 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>709,-54.5,711,-54.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>709 2</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>709,-62.5,711,-62.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>709 2</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>709,-70,711,-70</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>709 2</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>730,-58,730,-47</points>
<intersection>-58 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>730,-58,743,-58</points>
<connection>
<GID>84</GID>
<name>IN_3</name></connection>
<intersection>730 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>717,-47,730,-47</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>730 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>726,-59,743,-59</points>
<connection>
<GID>84</GID>
<name>IN_2</name></connection>
<intersection>726 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>726,-59,726,-55.5</points>
<intersection>-59 1</intersection>
<intersection>-55.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>717,-55.5,726,-55.5</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<intersection>726 3</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>730,-63.5,730,-60</points>
<intersection>-63.5 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>730,-60,743,-60</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>730 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>717,-63.5,730,-63.5</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>730 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>731,-71,731,-61</points>
<intersection>-71 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>731,-61,743,-61</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>731 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>717,-71,731,-71</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>731 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>607.695,274.549,1136.28,13.2789</PageViewport>
<gate>
<ID>36</ID>
<type>DD_KEYPAD_HEX</type>
<position>637.5,178.5</position>
<output>
<ID>OUT_0</ID>115 </output>
<output>
<ID>OUT_1</ID>114 </output>
<output>
<ID>OUT_2</ID>41 </output>
<output>
<ID>OUT_3</ID>38 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>51</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>720,178.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>114 </input>
<input>
<ID>IN_2</ID>41 </input>
<input>
<ID>IN_3</ID>38 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 15</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_TOGGLE</type>
<position>239.5,313</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>679.5,180.5,679.5,181.5</points>
<intersection>180.5 1</intersection>
<intersection>181.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>679.5,180.5,717,180.5</points>
<connection>
<GID>51</GID>
<name>IN_3</name></connection>
<intersection>679.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>642.5,181.5,679.5,181.5</points>
<connection>
<GID>36</GID>
<name>OUT_3</name></connection>
<intersection>679.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>642.5,179.5,717,179.5</points>
<connection>
<GID>51</GID>
<name>IN_2</name></connection>
<connection>
<GID>36</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>679.5,177.5,679.5,178.5</points>
<intersection>177.5 2</intersection>
<intersection>178.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>679.5,178.5,717,178.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>679.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>642.5,177.5,679.5,177.5</points>
<connection>
<GID>36</GID>
<name>OUT_1</name></connection>
<intersection>679.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>679.5,175.5,679.5,176</points>
<intersection>175.5 2</intersection>
<intersection>176 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>679.5,176,717,176</points>
<intersection>679.5 0</intersection>
<intersection>717 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>642.5,175.5,679.5,175.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>679.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>717,176,717,177.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>176 1</intersection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>-17.2648,1168.58,1206.74,563.581</PageViewport></page 3>
<page 4>
<PageViewport>-17.2648,1168.58,1206.74,563.581</PageViewport></page 4>
<page 5>
<PageViewport>-17.2648,1168.58,1206.74,563.581</PageViewport></page 5>
<page 6>
<PageViewport>-17.2648,1168.58,1206.74,563.581</PageViewport></page 6>
<page 7>
<PageViewport>-17.2648,1168.58,1206.74,563.581</PageViewport></page 7>
<page 8>
<PageViewport>-17.2648,1168.58,1206.74,563.581</PageViewport></page 8>
<page 9>
<PageViewport>-17.2648,1168.58,1206.74,563.581</PageViewport></page 9></circuit>
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>490.703,22.9378,877.985,-168.488</PageViewport>
<gate>
<ID>193</ID>
<type>AA_INVERTER</type>
<position>593.5,-102.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1</ID>
<type>AA_AND4</type>
<position>664,17.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>5 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>195</ID>
<type>AA_INVERTER</type>
<position>591.5,-106.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_FULLADDER_1BIT</type>
<position>584.5,-38</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_B_0</ID>9 </input>
<output>
<ID>OUT_0</ID>14 </output>
<input>
<ID>carry_in</ID>10 </input>
<output>
<ID>carry_out</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_FULLADDER_1BIT</type>
<position>567.5,-38</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_B_0</ID>8 </input>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>carry_in</ID>7 </input>
<output>
<ID>carry_out</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_INVERTER</type>
<position>591.5,-112</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5</ID>
<type>AI_XOR2</type>
<position>566.5,-29</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR2</type>
<position>578.5,-29</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AI_INVERTER_4BIT</type>
<position>658,27.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>1 </input>
<output>
<ID>OUT_0</ID>15 </output>
<output>
<ID>OUT_1</ID>16 </output>
<output>
<ID>OUT_2</ID>23 </output>
<output>
<ID>OUT_3</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>201</ID>
<type>AO_XNOR2</type>
<position>609.5,-121</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>561.5,23.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>561.5,20.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>203</ID>
<type>AO_XNOR2</type>
<position>609.5,-126</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>561.5,17</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>561.5,13.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_AND2</type>
<position>637,-129</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>555.5,24</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>555.5,21</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_AND3</type>
<position>609,-134</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>97 </input>
<input>
<ID>IN_2</ID>98 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>555.5,17.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>555.5,14</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_AND3</type>
<position>609,-141</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>1 </input>
<input>
<ID>IN_2</ID>99 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>707.5,47.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>707,43</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_AND2</type>
<position>609,-147</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>561.5,-11</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>213</ID>
<type>AE_OR3</type>
<position>638,-139.5</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>110 </input>
<input>
<ID>IN_2</ID>111 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_OR4</type>
<position>660.5,6.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>5 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>21</ID>
<type>AI_XOR4</type>
<position>662,-4</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>5 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_INVERTER</type>
<position>671.5,12.5</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_INVERTER</type>
<position>674,4</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_INVERTER</type>
<position>591,-134</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_INVERTER</type>
<position>673,-8.5</position>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AI_MUX_8x1</type>
<position>691.5,25.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>19 </input>
<input>
<ID>IN_3</ID>11 </input>
<input>
<ID>IN_4</ID>15 </input>
<input>
<ID>IN_5</ID>16 </input>
<input>
<ID>IN_6</ID>23 </input>
<input>
<ID>IN_7</ID>17 </input>
<output>
<ID>OUT</ID>24 </output>
<input>
<ID>SEL_0</ID>13 </input>
<input>
<ID>SEL_1</ID>12 </input>
<input>
<ID>SEL_2</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>219</ID>
<type>AA_INVERTER</type>
<position>597,-136</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_MUX_2x1</type>
<position>717.5,24.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>27 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>767.5,24.5</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AA_INVERTER</type>
<position>596,-143</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>694.5,47.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>699,47.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AA_INVERTER</type>
<position>591,-148</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>703.5,47.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>695.5,43</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>699.5,43</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>703.5,43</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>768.5,-113.5</position>
<gparam>LABEL_TEXT A  B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>608.5,-49</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>608.5,-54</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>768.5,-124.5</position>
<gparam>LABEL_TEXT A = B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_AND2</type>
<position>608.5,-59</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>608.5,-64</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>769,-135.5</position>
<gparam>LABEL_TEXT A > B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AI_XOR2</type>
<position>646.5,-52.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_AND2</type>
<position>643.5,-57</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AI_MUX_8x1</type>
<position>703.5,-22</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>107 </input>
<input>
<ID>IN_2</ID>101 </input>
<input>
<ID>IN_3</ID>22 </input>
<input>
<ID>IN_4</ID>7 </input>
<input>
<ID>IN_5</ID>14 </input>
<input>
<ID>IN_6</ID>4 </input>
<input>
<ID>IN_7</ID>18 </input>
<output>
<ID>OUT</ID>36 </output>
<input>
<ID>SEL_0</ID>13 </input>
<input>
<ID>SEL_1</ID>12 </input>
<input>
<ID>SEL_2</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>47</ID>
<type>AI_XOR2</type>
<position>655.5,-59.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_AND2</type>
<position>656.5,-66.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>767.5,3.5</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>646,-107.5</position>
<gparam>LABEL_TEXT COMPARATOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>768,-21</position>
<gparam>LABEL_TEXT MUL</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>768,-44.5</position>
<gparam>LABEL_TEXT DIV</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>537,18.5</position>
<gparam>LABEL_TEXT INPUTS</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>682.5,38.5</position>
<gparam>LABEL_TEXT SELECT LINES</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>768.5,-118.5</position>
<input>
<ID>N_in0</ID>101 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>768,-29.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<input>
<ID>IN_2</ID>34 </input>
<input>
<ID>IN_3</ID>35 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>766.5,29</position>
<gparam>LABEL_TEXT Output</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>GA_LED</type>
<position>768.5,-129</position>
<input>
<ID>N_in0</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>765,7.5</position>
<gparam>LABEL_TEXT Int. C/ B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>553,-10.5</position>
<gparam>LABEL_TEXT Key A/ S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>768.5,-139.5</position>
<input>
<ID>N_in0</ID>108 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_AND3</type>
<position>677,-71.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>49 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_INVERTER</type>
<position>656.5,-73.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_OR2</type>
<position>675,-79</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_AND3</type>
<position>690,-81</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>1 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND3</type>
<position>670.5,-87</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>51 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_INVERTER</type>
<position>657.5,-89</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR3</type>
<position>714.5,-80</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>54 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND3</type>
<position>668.5,-94</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>56 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_INVERTER</type>
<position>646,-96</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>123</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>768,-52.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>57 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>612.5,-28.5</position>
<gparam>LABEL_TEXT ADDER/ SUB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>708,-75</position>
<gparam>LABEL_TEXT MULTIPLIER</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AA_LABEL</type>
<position>679,-90.5</position>
<gparam>LABEL_TEXT DIVIDER</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_AND3</type>
<position>609.5,-100.5</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_2</ID>2 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_AND2</type>
<position>609.5,-107.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_AND3</type>
<position>609.5,-114</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>2 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>189</ID>
<type>AE_OR3</type>
<position>637.5,-118.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>86 </input>
<input>
<ID>IN_2</ID>87 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_INVERTER</type>
<position>590,-98.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>624,-12.5,624,23.5</points>
<intersection>-12.5 28</intersection>
<intersection>-1 26</intersection>
<intersection>9.5 14</intersection>
<intersection>21.5 4</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>563.5,23.5,656,23.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>624 0</intersection>
<intersection>656 50</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>624,21.5,659.5,21.5</points>
<intersection>624 0</intersection>
<intersection>659.5 51</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>624,9.5,657.5,9.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>624 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>624,-1,659,-1</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>624 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>601,-12.5,624,-12.5</points>
<intersection>601 30</intersection>
<intersection>624 0</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>601,-48,601,-12.5</points>
<intersection>-48 31</intersection>
<intersection>-35 32</intersection>
<intersection>-12.5 28</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>593.5,-48,605.5,-48</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>593.5 33</intersection>
<intersection>601 30</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>585.5,-35,601,-35</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>601 30</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>593.5,-58,593.5,-48</points>
<intersection>-58 34</intersection>
<intersection>-48 31</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>572.5,-58,605.5,-58</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>572.5 36</intersection>
<intersection>593.5 33</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>572.5,-69.5,572.5,-58</points>
<intersection>-69.5 37</intersection>
<intersection>-58 34</intersection></vsegment>
<hsegment>
<ID>37</ID>
<points>561,-69.5,674,-69.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>561 38</intersection>
<intersection>572.5 36</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>561,-83,561,-69.5</points>
<intersection>-83 39</intersection>
<intersection>-69.5 37</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>561,-83,687,-83</points>
<connection>
<GID>115</GID>
<name>IN_2</name></connection>
<intersection>561 38</intersection>
<intersection>567.5 40</intersection></hsegment>
<vsegment>
<ID>40</ID>
<points>567.5,-102.5,567.5,-83</points>
<intersection>-102.5 41</intersection>
<intersection>-83 39</intersection></vsegment>
<hsegment>
<ID>41</ID>
<points>559,-102.5,590.5,-102.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>559 42</intersection>
<intersection>567.5 40</intersection></hsegment>
<vsegment>
<ID>42</ID>
<points>559,-141,559,-102.5</points>
<intersection>-141 49</intersection>
<intersection>-132 47</intersection>
<intersection>-125 45</intersection>
<intersection>-112 43</intersection>
<intersection>-102.5 41</intersection></vsegment>
<hsegment>
<ID>43</ID>
<points>559,-112,588.5,-112</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>559 42</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>559,-125,606.5,-125</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>559 42</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>559,-132,606,-132</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>559 42</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>559,-141,606,-141</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>559 42</intersection></hsegment>
<vsegment>
<ID>50</ID>
<points>656,23.5,656,29</points>
<connection>
<GID>7</GID>
<name>IN_3</name></connection>
<intersection>23.5 1</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>659.5,20.5,659.5,21.5</points>
<intersection>20.5 52</intersection>
<intersection>21.5 4</intersection></vsegment>
<hsegment>
<ID>52</ID>
<points>659.5,20.5,661,20.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>659.5 51</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>627,-19,627,28</points>
<intersection>-19 26</intersection>
<intersection>-3 23</intersection>
<intersection>7.5 14</intersection>
<intersection>20.5 2</intersection>
<intersection>28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>627,28,656,28</points>
<connection>
<GID>7</GID>
<name>IN_2</name></connection>
<intersection>627 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>563.5,20.5,654,20.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>627 0</intersection>
<intersection>654 56</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>627,7.5,657.5,7.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>627 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>627,-3,659,-3</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>627 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>577.5,-19,627,-19</points>
<intersection>577.5 27</intersection>
<intersection>598 33</intersection>
<intersection>627 0</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>577.5,-26,577.5,-19</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-19 26</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>598,-50,598,-19</points>
<intersection>-50 34</intersection>
<intersection>-19 26</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>598,-50,605.5,-50</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>598 33</intersection>
<intersection>601 35</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>601,-55,601,-50</points>
<intersection>-55 36</intersection>
<intersection>-50 34</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>562.5,-55,605.5,-55</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>562.5 38</intersection>
<intersection>601 35</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>562.5,-71.5,562.5,-55</points>
<intersection>-71.5 39</intersection>
<intersection>-55 36</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>562.5,-71.5,674,-71.5</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>562.5 38</intersection>
<intersection>636.5 40</intersection></hsegment>
<vsegment>
<ID>40</ID>
<points>636.5,-78,636.5,-71.5</points>
<intersection>-78 41</intersection>
<intersection>-71.5 39</intersection></vsegment>
<hsegment>
<ID>41</ID>
<points>615.5,-78,672,-78</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>615.5 42</intersection>
<intersection>636.5 40</intersection></hsegment>
<vsegment>
<ID>42</ID>
<points>615.5,-89,615.5,-78</points>
<intersection>-89 43</intersection>
<intersection>-78 41</intersection></vsegment>
<hsegment>
<ID>43</ID>
<points>563,-89,654.5,-89</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>563 44</intersection>
<intersection>615.5 42</intersection></hsegment>
<vsegment>
<ID>44</ID>
<points>563,-94,563,-89</points>
<intersection>-94 45</intersection>
<intersection>-89 43</intersection></vsegment>
<hsegment>
<ID>45</ID>
<points>563,-94,665.5,-94</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>563 44</intersection>
<intersection>573.5 46</intersection></hsegment>
<vsegment>
<ID>46</ID>
<points>573.5,-104.5,573.5,-94</points>
<intersection>-104.5 47</intersection>
<intersection>-94 45</intersection></vsegment>
<hsegment>
<ID>47</ID>
<points>564.5,-104.5,597.5,-104.5</points>
<intersection>564.5 48</intersection>
<intersection>573.5 46</intersection>
<intersection>597.5 57</intersection></hsegment>
<vsegment>
<ID>48</ID>
<points>564.5,-143,564.5,-104.5</points>
<intersection>-143 55</intersection>
<intersection>-136 53</intersection>
<intersection>-127 51</intersection>
<intersection>-116 49</intersection>
<intersection>-104.5 47</intersection></vsegment>
<hsegment>
<ID>49</ID>
<points>564.5,-116,606.5,-116</points>
<connection>
<GID>187</GID>
<name>IN_2</name></connection>
<intersection>564.5 48</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>564.5,-127,606.5,-127</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>564.5 48</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>564.5,-136,594,-136</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>564.5 48</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>564.5,-143,593,-143</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>564.5 48</intersection></hsegment>
<vsegment>
<ID>56</ID>
<points>654,18.5,654,20.5</points>
<intersection>18.5 59</intersection>
<intersection>20.5 2</intersection></vsegment>
<vsegment>
<ID>57</ID>
<points>597.5,-104.5,597.5,-102.5</points>
<intersection>-104.5 47</intersection>
<intersection>-102.5 58</intersection></vsegment>
<hsegment>
<ID>58</ID>
<points>597.5,-102.5,606.5,-102.5</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>597.5 57</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>654,18.5,661,18.5</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>654 56</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>688,-19.5,688,-8.5</points>
<intersection>-19.5 3</intersection>
<intersection>-8.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>688,-19.5,700.5,-19.5</points>
<connection>
<GID>46</GID>
<name>IN_6</name></connection>
<intersection>688 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>676,-8.5,688,-8.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>688 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>630.5,-16.5,630.5,27</points>
<intersection>-16.5 28</intersection>
<intersection>-5 26</intersection>
<intersection>5.5 18</intersection>
<intersection>17 15</intersection>
<intersection>27 22</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>563.5,17,661,17</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>630.5 0</intersection>
<intersection>661 35</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>630.5,5.5,657.5,5.5</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>630.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>630.5,27,656,27</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>630.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>630.5,-5,659,-5</points>
<connection>
<GID>21</GID>
<name>IN_2</name></connection>
<intersection>630.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>559,-16.5,630.5,-16.5</points>
<intersection>559 30</intersection>
<intersection>630.5 0</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>559,-98.5,559,-16.5</points>
<intersection>-98.5 44</intersection>
<intersection>-85 40</intersection>
<intersection>-81 38</intersection>
<intersection>-53 31</intersection>
<intersection>-35 32</intersection>
<intersection>-16.5 28</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>559,-53,605.5,-53</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>559 30</intersection>
<intersection>582 33</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>559,-35,568.5,-35</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>559 30</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>582,-63,582,-53</points>
<intersection>-63 34</intersection>
<intersection>-53 31</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>566,-63,605.5,-63</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>566 37</intersection>
<intersection>582 33</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>661,16.5,661,17</points>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>17 15</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>566,-81,566,-63</points>
<intersection>-81 38</intersection>
<intersection>-63 34</intersection></vsegment>
<hsegment>
<ID>38</ID>
<points>559,-81,687,-81</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>559 30</intersection>
<intersection>566 37</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>559,-85,667.5,-85</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>559 30</intersection>
<intersection>614 41</intersection></hsegment>
<vsegment>
<ID>41</ID>
<points>614,-92,614,-85</points>
<intersection>-92 42</intersection>
<intersection>-85 40</intersection></vsegment>
<hsegment>
<ID>42</ID>
<points>614,-92,665.5,-92</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>614 41</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>559,-98.5,587,-98.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>559 30</intersection>
<intersection>583.5 45</intersection></hsegment>
<vsegment>
<ID>45</ID>
<points>583.5,-106.5,583.5,-98.5</points>
<intersection>-106.5 46</intersection>
<intersection>-98.5 44</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>567,-106.5,588.5,-106.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>567 47</intersection>
<intersection>583.5 45</intersection></hsegment>
<vsegment>
<ID>47</ID>
<points>567,-146,567,-106.5</points>
<intersection>-146 52</intersection>
<intersection>-139 50</intersection>
<intersection>-120 48</intersection>
<intersection>-106.5 46</intersection></vsegment>
<hsegment>
<ID>48</ID>
<points>567,-120,606.5,-120</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>567 47</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>567,-139,606,-139</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>567 47</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>567,-146,606,-146</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>567 47</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>634.5,-7,634.5,26</points>
<intersection>-7 4</intersection>
<intersection>3.5 7</intersection>
<intersection>14.5 6</intersection>
<intersection>26 24</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>620.5,-7,659,-7</points>
<connection>
<GID>21</GID>
<name>IN_3</name></connection>
<intersection>620.5 12</intersection>
<intersection>634.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>634.5,14.5,661,14.5</points>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>634.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>634.5,3.5,657.5,3.5</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<intersection>634.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>620.5,-16.5,620.5,13.5</points>
<intersection>-16.5 21</intersection>
<intersection>-7 4</intersection>
<intersection>13.5 27</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>565.5,-16.5,620.5,-16.5</points>
<intersection>565.5 22</intersection>
<intersection>600 28</intersection>
<intersection>620.5 12</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>565.5,-26,565.5,-16.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>-16.5 21</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>634.5,26,656,26</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>634.5 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>563.5,13.5,620.5,13.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>620.5 12</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>600,-65,600,-16.5</points>
<intersection>-65 30</intersection>
<intersection>-60 29</intersection>
<intersection>-16.5 21</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>600,-60,605.5,-60</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>600 28</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>588,-65,605.5,-65</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>588 31</intersection>
<intersection>600 28</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>588,-73.5,588,-65</points>
<intersection>-73.5 32</intersection>
<intersection>-65 30</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>588,-73.5,653.5,-73.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>588 31</intersection>
<intersection>648 33</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>648,-80,648,-73.5</points>
<intersection>-80 34</intersection>
<intersection>-73.5 32</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>624.5,-80,672,-80</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>624.5 35</intersection>
<intersection>648 33</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>624.5,-87,624.5,-80</points>
<intersection>-87 36</intersection>
<intersection>-80 34</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>561,-87,667.5,-87</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>561 37</intersection>
<intersection>624.5 35</intersection></hsegment>
<vsegment>
<ID>37</ID>
<points>561,-148,561,-87</points>
<intersection>-148 48</intersection>
<intersection>-134 46</intersection>
<intersection>-122 44</intersection>
<intersection>-114 42</intersection>
<intersection>-108.5 40</intersection>
<intersection>-96 38</intersection>
<intersection>-87 36</intersection></vsegment>
<hsegment>
<ID>38</ID>
<points>561,-96,643,-96</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>561 37</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>561,-108.5,606.5,-108.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>561 37</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>561,-114,606.5,-114</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>561 37</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>561,-122,606.5,-122</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>561 37</intersection>
<intersection>584.5 45</intersection></hsegment>
<vsegment>
<ID>45</ID>
<points>584.5,-134,584.5,-122</points>
<intersection>-134 46</intersection>
<intersection>-122 44</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>561,-134,588,-134</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>561 37</intersection>
<intersection>584.5 45</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>561,-148,588,-148</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>561 37</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>571.5,-43,693.5,-43</points>
<intersection>571.5 14</intersection>
<intersection>580.5 13</intersection>
<intersection>693.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>693.5,-43,693.5,-21.5</points>
<intersection>-43 6</intersection>
<intersection>-21.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>693.5,-21.5,700.5,-21.5</points>
<connection>
<GID>46</GID>
<name>IN_4</name></connection>
<intersection>693.5 9</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>580.5,-43,580.5,-38</points>
<connection>
<GID>2</GID>
<name>carry_out</name></connection>
<intersection>-43 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>571.5,-43,571.5,-38</points>
<connection>
<GID>3</GID>
<name>carry_in</name></connection>
<intersection>-43 6</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>566.5,-35,566.5,-32</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<connection>
<GID>3</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583.5,-35,583.5,-32</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<intersection>-32 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>578.5,-32,583.5,-32</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>583.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593.5,-38,593.5,-11</points>
<intersection>-38 3</intersection>
<intersection>-24.5 4</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>563.5,-11,593.5,-11</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>567.5 2</intersection>
<intersection>593.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>567.5,-26,567.5,-11</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>588.5,-38,593.5,-38</points>
<connection>
<GID>2</GID>
<name>carry_in</name></connection>
<intersection>593.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>579.5,-24.5,593.5,-24.5</points>
<intersection>579.5 5</intersection>
<intersection>593.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>579.5,-26,579.5,-24.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-24.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>667,17.5,677,17.5</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<intersection>667 4</intersection>
<intersection>677 13</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>667,12.5,667,17.5</points>
<intersection>12.5 5</intersection>
<intersection>17.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>667,12.5,668.5,12.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>667 4</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>677,17.5,677,25</points>
<intersection>17.5 1</intersection>
<intersection>25 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>677,25,688.5,25</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>677 13</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>703.5,-16.5,703.5,35</points>
<connection>
<GID>46</GID>
<name>SEL_1</name></connection>
<intersection>32 6</intersection>
<intersection>35 10</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>691.5,32,703.5,32</points>
<intersection>691.5 11</intersection>
<intersection>703.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>699.5,35,703.5,35</points>
<intersection>699.5 12</intersection>
<intersection>703.5 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>691.5,31,691.5,32</points>
<connection>
<GID>25</GID>
<name>SEL_1</name></connection>
<intersection>32 6</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>699.5,35,699.5,41</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>35 10</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>704.5,-16.5,704.5,41</points>
<connection>
<GID>46</GID>
<name>SEL_0</name></connection>
<intersection>31.5 15</intersection>
<intersection>41 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>703.5,41,704.5,41</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>704.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>692.5,31.5,704.5,31.5</points>
<intersection>692.5 16</intersection>
<intersection>704.5 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>692.5,31,692.5,31.5</points>
<connection>
<GID>25</GID>
<name>SEL_0</name></connection>
<intersection>31.5 15</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584.5,-41,584.5,-20.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>584.5,-20.5,700.5,-20.5</points>
<connection>
<GID>46</GID>
<name>IN_5</name></connection>
<intersection>584.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>660,26,688.5,26</points>
<connection>
<GID>25</GID>
<name>IN_4</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>660,27,688.5,27</points>
<connection>
<GID>25</GID>
<name>IN_5</name></connection>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>660,29,688.5,29</points>
<connection>
<GID>25</GID>
<name>IN_7</name></connection>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>666,-4,670,-4</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>670 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>670,-18.5,670,-4</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-18.5 11</intersection>
<intersection>-4 7</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>670,-18.5,700.5,-18.5</points>
<connection>
<GID>46</GID>
<name>IN_7</name></connection>
<intersection>670 9</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>679,24,688.5,24</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>679 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>679,12.5,679,24</points>
<intersection>12.5 5</intersection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>674.5,12.5,679,12.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>679 4</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>664.5,6.5,681.5,6.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>664.5 3</intersection>
<intersection>681.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>664.5,4,664.5,6.5</points>
<intersection>4 4</intersection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>664.5,4,671,4</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>664.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>681.5,6.5,681.5,23</points>
<intersection>6.5 1</intersection>
<intersection>23 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>681.5,23,688.5,23</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>681.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>684.5,4,684.5,22</points>
<intersection>4 3</intersection>
<intersection>22 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>677,4,684.5,4</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>684.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>684.5,22,688.5,22</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>684.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>569.5,-41,569.5,-22.5</points>
<intersection>-41 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>569.5,-22.5,700.5,-22.5</points>
<connection>
<GID>46</GID>
<name>IN_3</name></connection>
<intersection>569.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>567.5,-41,569.5,-41</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>569.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>660,28,688.5,28</points>
<connection>
<GID>25</GID>
<name>IN_6</name></connection>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>694.5,25.5,715.5,25.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<connection>
<GID>25</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>707,27,707,41</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>707,27,717.5,27</points>
<connection>
<GID>26</GID>
<name>SEL_0</name></connection>
<intersection>707 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>702.5,-16.5,702.5,34</points>
<connection>
<GID>46</GID>
<name>SEL_2</name></connection>
<intersection>33 6</intersection>
<intersection>34 10</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>690.5,33,702.5,33</points>
<intersection>690.5 13</intersection>
<intersection>702.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>695.5,34,702.5,34</points>
<intersection>695.5 11</intersection>
<intersection>702.5 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>695.5,34,695.5,41</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>34 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>690.5,31,690.5,33</points>
<connection>
<GID>25</GID>
<name>SEL_2</name></connection>
<intersection>33 6</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>719.5,24.5,766.5,24.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>27</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>623,-54,623,-51.5</points>
<intersection>-54 2</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>623,-51.5,643.5,-51.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>623 0</intersection>
<intersection>635.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>611.5,-54,623,-54</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>623 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>635.5,-56,635.5,-51.5</points>
<intersection>-56 4</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>635.5,-56,640.5,-56</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>635.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>624.5,-59,624.5,-53.5</points>
<intersection>-59 2</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>624.5,-53.5,643.5,-53.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>624.5 0</intersection>
<intersection>631.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>611.5,-59,624.5,-59</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>624.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>631.5,-58,631.5,-53.5</points>
<intersection>-58 4</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>631.5,-58,640.5,-58</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>631.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>647.5,-58.5,647.5,-57</points>
<intersection>-58.5 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>647.5,-58.5,652.5,-58.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>647.5 0</intersection>
<intersection>649.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>646.5,-57,647.5,-57</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>647.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>649.5,-65.5,649.5,-58.5</points>
<intersection>-65.5 4</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>649.5,-65.5,653.5,-65.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>649.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>630,-64,630,-60.5</points>
<intersection>-64 2</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>630,-60.5,652.5,-60.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>630 0</intersection>
<intersection>646.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>611.5,-64,630,-64</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>630 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>646.5,-67.5,646.5,-60.5</points>
<intersection>-67.5 4</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>646.5,-67.5,653.5,-67.5</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>646.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>673,-56,673,-49</points>
<intersection>-56 1</intersection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>673,-56,736,-56</points>
<intersection>673 0</intersection>
<intersection>736 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>611.5,-49,673,-49</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<intersection>673 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>736,-56,736,-30.5</points>
<intersection>-56 1</intersection>
<intersection>-30.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>736,-30.5,765,-30.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>736 5</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>690,-62,690,-52.5</points>
<intersection>-62 1</intersection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>690,-62,734.5,-62</points>
<intersection>690 0</intersection>
<intersection>734.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>649.5,-52.5,690,-52.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>690 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>734.5,-62,734.5,-29.5</points>
<intersection>-62 1</intersection>
<intersection>-29.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>734.5,-29.5,765,-29.5</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>734.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>698,-69,698,-59.5</points>
<intersection>-69 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>698,-69,733.5,-69</points>
<intersection>698 0</intersection>
<intersection>733.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>658.5,-59.5,698,-59.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>698 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>733.5,-69,733.5,-28.5</points>
<intersection>-69 1</intersection>
<intersection>-28.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>733.5,-28.5,765,-28.5</points>
<connection>
<GID>63</GID>
<name>IN_2</name></connection>
<intersection>733.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>659.5,-66.5,732.5,-66.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>732.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>732.5,-66.5,732.5,-27.5</points>
<intersection>-66.5 1</intersection>
<intersection>-27.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>732.5,-27.5,765,-27.5</points>
<connection>
<GID>63</GID>
<name>IN_3</name></connection>
<intersection>732.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>711,-22,711,23.5</points>
<intersection>-22 3</intersection>
<intersection>23.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>706.5,-22,711,-22</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>711 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>711,23.5,715.5,23.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>711 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>563.5,-46,729.5,-46</points>
<intersection>563.5 4</intersection>
<intersection>729.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>729.5,-46,729.5,3.5</points>
<intersection>-46 1</intersection>
<intersection>3.5 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>563.5,-46,563.5,-38</points>
<connection>
<GID>3</GID>
<name>carry_out</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>729.5,3.5,766.5,3.5</points>
<connection>
<GID>50</GID>
<name>N_in0</name></connection>
<intersection>729.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>659.5,-73.5,674,-73.5</points>
<connection>
<GID>112</GID>
<name>IN_2</name></connection>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>678,-79,687,-79</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<connection>
<GID>115</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>660.5,-89,667.5,-89</points>
<connection>
<GID>116</GID>
<name>IN_2</name></connection>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>693,-81,708.5,-81</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>708.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>708.5,-81,708.5,-80</points>
<intersection>-81 1</intersection>
<intersection>-80 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>708.5,-80,711.5,-80</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>708.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>692.5,-78,692.5,-71.5</points>
<intersection>-78 1</intersection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>692.5,-78,711.5,-78</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>692.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>680,-71.5,692.5,-71.5</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>692.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673.5,-87,708.5,-87</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>708.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>708.5,-87,708.5,-82</points>
<intersection>-87 1</intersection>
<intersection>-82 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>708.5,-82,711.5,-82</points>
<connection>
<GID>118</GID>
<name>IN_2</name></connection>
<intersection>708.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>720,-99,720,-80</points>
<intersection>-99 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>720,-99,758,-99</points>
<intersection>720 0</intersection>
<intersection>758 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>717.5,-80,720,-80</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>720 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>758,-99,758,-53.5</points>
<intersection>-99 1</intersection>
<intersection>-53.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>758,-53.5,765,-53.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>758 7</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649,-96,665.5,-96</points>
<connection>
<GID>120</GID>
<name>IN_2</name></connection>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>699.5,-104.5,699.5,-94</points>
<intersection>-104.5 1</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>699.5,-104.5,760.5,-104.5</points>
<intersection>699.5 0</intersection>
<intersection>760.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>671.5,-94,699.5,-94</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>699.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>760.5,-104.5,760.5,-52.5</points>
<intersection>-104.5 1</intersection>
<intersection>-52.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>760.5,-52.5,765,-52.5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>760.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>631.5,-116.5,631.5,-100.5</points>
<intersection>-116.5 1</intersection>
<intersection>-100.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>631.5,-116.5,634.5,-116.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>631.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>612.5,-100.5,631.5,-100.5</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<intersection>631.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612.5,-107.5,629.5,-107.5</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>629.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>629.5,-118.5,629.5,-107.5</points>
<intersection>-118.5 3</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>629.5,-118.5,634.5,-118.5</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<intersection>629.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>622.5,-120.5,622.5,-114</points>
<intersection>-120.5 2</intersection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>612.5,-114,622.5,-114</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<intersection>622.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>622.5,-120.5,634.5,-120.5</points>
<connection>
<GID>189</GID>
<name>IN_2</name></connection>
<intersection>622.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593,-98.5,606.5,-98.5</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<connection>
<GID>183</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>597,-100.5,606.5,-100.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>597 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>597,-102.5,597,-100.5</points>
<intersection>-102.5 9</intersection>
<intersection>-100.5 0</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>596.5,-102.5,597,-102.5</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<intersection>597 8</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>594.5,-106.5,606.5,-106.5</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<connection>
<GID>185</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>594.5,-112,606.5,-112</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>594,-134,606,-134</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600,-136,606,-136</points>
<connection>
<GID>207</GID>
<name>IN_2</name></connection>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>599,-143,606,-143</points>
<connection>
<GID>209</GID>
<name>IN_2</name></connection>
<connection>
<GID>221</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>594,-148,606,-148</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>640.5,-118.5,767.5,-118.5</points>
<connection>
<GID>189</GID>
<name>OUT</name></connection>
<connection>
<GID>62</GID>
<name>N_in0</name></connection>
<intersection>696.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>696.5,-118.5,696.5,-23.5</points>
<intersection>-118.5 1</intersection>
<intersection>-23.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>696.5,-23.5,700.5,-23.5</points>
<connection>
<GID>46</GID>
<name>IN_2</name></connection>
<intersection>696.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>623.5,-128,623.5,-121</points>
<intersection>-128 1</intersection>
<intersection>-121 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>623.5,-128,634,-128</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>623.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>612.5,-121,623.5,-121</points>
<connection>
<GID>201</GID>
<name>OUT</name></connection>
<intersection>623.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>614,-130,634,-130</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>614 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>614,-130,614,-126</points>
<intersection>-130 1</intersection>
<intersection>-126 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>612.5,-126,614,-126</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>614 3</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>640,-129,767.5,-129</points>
<connection>
<GID>205</GID>
<name>OUT</name></connection>
<connection>
<GID>66</GID>
<name>N_in0</name></connection>
<intersection>695.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>695.5,-129,695.5,-24.5</points>
<intersection>-129 1</intersection>
<intersection>-24.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>695.5,-24.5,700.5,-24.5</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>695.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>641,-139.5,767.5,-139.5</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<connection>
<GID>70</GID>
<name>N_in0</name></connection>
<intersection>694.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>694.5,-139.5,694.5,-25.5</points>
<intersection>-139.5 1</intersection>
<intersection>-25.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>694.5,-25.5,700.5,-25.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>694.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612,-137.5,635,-137.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>612 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>612,-137.5,612,-134</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<intersection>-137.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>623,-141,623,-139.5</points>
<intersection>-141 2</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>623,-139.5,635,-139.5</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>623 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>612,-141,623,-141</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<intersection>623 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>624,-147,624,-141.5</points>
<intersection>-147 2</intersection>
<intersection>-141.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>624,-141.5,635,-141.5</points>
<connection>
<GID>213</GID>
<name>IN_2</name></connection>
<intersection>624 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>612,-147,624,-147</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>624 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>119.143,21.134,726.341,-278.992</PageViewport>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>184.5,-45.5</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>177,-45.5</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_TOGGLE</type>
<position>169.5,-45.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_TOGGLE</type>
<position>162,-45.5</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>161,-42</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>169.5,-41.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>177,-41.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>184.5,-41.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_AND3</type>
<position>220,-57</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>69 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_INVERTER</type>
<position>205.5,-62</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_INVERTER</type>
<position>199,-64.5</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_AND2</type>
<position>213,-71.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_AND3</type>
<position>213,-78.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>71 </input>
<input>
<ID>IN_2</ID>69 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>141</ID>
<type>AE_OR3</type>
<position>237,-70.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>60 </input>
<input>
<ID>IN_2</ID>61 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_OR2</type>
<position>60.5,-57</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND2</type>
<position>231,-88</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_AND3</type>
<position>213,-107.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>74 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_AND2</type>
<position>213,-114</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AE_OR3</type>
<position>233.5,-107</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>65 </input>
<input>
<ID>IN_2</ID>66 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_INVERTER</type>
<position>204,-72.5</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_INVERTER</type>
<position>207,-76.5</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_INVERTER</type>
<position>206.5,-98</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_INVERTER</type>
<position>207,-109.5</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_INVERTER</type>
<position>207,-115</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>252,-70</position>
<input>
<ID>N_in0</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>GA_LED</type>
<position>252,-87.5</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>GA_LED</type>
<position>252.5,-104.5</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AO_XNOR2</type>
<position>202.5,-85.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>71 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AO_XNOR2</type>
<position>202.5,-91.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_AND3</type>
<position>217.5,-98.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>84 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_INVERTER</type>
<position>209,-102</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206,-64.5,206,-57</points>
<intersection>-64.5 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206,-57,217,-57</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>206 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>202,-64.5,206,-64.5</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<intersection>206 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-68.5,225,-57</points>
<intersection>-68.5 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,-68.5,234,-68.5</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,-57,225,-57</points>
<connection>
<GID>131</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-71.5,225,-70.5</points>
<intersection>-71.5 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,-70.5,234,-70.5</points>
<connection>
<GID>141</GID>
<name>IN_1</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-71.5,225,-71.5</points>
<connection>
<GID>137</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-78.5,225,-72.5</points>
<intersection>-78.5 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,-72.5,234,-72.5</points>
<connection>
<GID>141</GID>
<name>IN_2</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-78.5,225,-78.5</points>
<connection>
<GID>139</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223,-107.5,223,-107</points>
<intersection>-107.5 2</intersection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223,-107,230.5,-107</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>223 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-107.5,223,-107.5</points>
<connection>
<GID>153</GID>
<name>OUT</name></connection>
<intersection>223 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223,-114,223,-109</points>
<intersection>-114 2</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223,-109,230.5,-109</points>
<connection>
<GID>157</GID>
<name>IN_2</name></connection>
<intersection>223 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-114,223,-114</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<intersection>223 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-62,177,-47.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,-62,202.5,-62</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>177 0</intersection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-72.5,192,-62</points>
<intersection>-72.5 3</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-72.5,201,-72.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>176 4</intersection>
<intersection>180.5 10</intersection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>176,-113,176,-72.5</points>
<intersection>-113 9</intersection>
<intersection>-105.5 7</intersection>
<intersection>-72.5 3</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>176,-105.5,210,-105.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>176 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>176,-113,210,-113</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>176 4</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>180.5,-84.5,180.5,-72.5</points>
<intersection>-84.5 11</intersection>
<intersection>-72.5 3</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>180.5,-84.5,199.5,-84.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>180.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-107.5,162,-47.5</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<intersection>-107.5 9</intersection>
<intersection>-98.5 7</intersection>
<intersection>-76.5 3</intersection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162,-64.5,196,-64.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>162,-76.5,204,-76.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>162,-98.5,164,-98.5</points>
<intersection>162 0</intersection>
<intersection>164 10</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>162,-107.5,210,-107.5</points>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<intersection>162 0</intersection>
<intersection>196 12</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>164,-98.5,164,-90.5</points>
<intersection>-98.5 7</intersection>
<intersection>-90.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>164,-90.5,199.5,-90.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>164 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>196,-107.5,196,-96.5</points>
<intersection>-107.5 9</intersection>
<intersection>-96.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>196,-96.5,214.5,-96.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>196 12</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-109.5,169.5,-47.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 9</intersection>
<intersection>-102.5 7</intersection>
<intersection>-80.5 3</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-59,217,-59</points>
<connection>
<GID>131</GID>
<name>IN_2</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>169.5,-80.5,210,-80.5</points>
<connection>
<GID>139</GID>
<name>IN_2</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>169.5,-102.5,193,-102.5</points>
<intersection>169.5 0</intersection>
<intersection>193 10</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>169.5,-109.5,204,-109.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection>
<intersection>201.5 12</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>193,-102.5,193,-92.5</points>
<intersection>-102.5 7</intersection>
<intersection>-92.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>193,-92.5,199.5,-92.5</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>193 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>201.5,-109.5,201.5,-102</points>
<intersection>-109.5 9</intersection>
<intersection>-102 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>201.5,-102,206,-102</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>201.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>207,-72.5,210,-72.5</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-115,184.5,-47.5</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>-115 9</intersection>
<intersection>-98 7</intersection>
<intersection>-78.5 3</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,-70.5,210,-70.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>184.5,-78.5,210,-78.5</points>
<connection>
<GID>139</GID>
<name>IN_1</name></connection>
<intersection>184.5 0</intersection>
<intersection>186.5 10</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>184.5,-98,203.5,-98</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>184.5,-115,204,-115</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>186.5,-86.5,186.5,-78.5</points>
<intersection>-86.5 11</intersection>
<intersection>-78.5 3</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>186.5,-86.5,199.5,-86.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>186.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-76.5,210,-76.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-109.5,210,-109.5</points>
<connection>
<GID>153</GID>
<name>IN_2</name></connection>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-115,210,-115</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-70.5,245.5,-70</points>
<intersection>-70.5 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245.5,-70,251,-70</points>
<connection>
<GID>169</GID>
<name>N_in0</name></connection>
<intersection>245.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>240,-70.5,245.5,-70.5</points>
<connection>
<GID>141</GID>
<name>OUT</name></connection>
<intersection>245.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242.5,-88,242.5,-87.5</points>
<intersection>-88 2</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242.5,-87.5,251,-87.5</points>
<connection>
<GID>171</GID>
<name>N_in0</name></connection>
<intersection>242.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234,-88,242.5,-88</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>242.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-107,244,-104.5</points>
<intersection>-107 2</intersection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,-104.5,251.5,-104.5</points>
<connection>
<GID>173</GID>
<name>N_in0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>236.5,-107,244,-107</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216.5,-87,216.5,-85.5</points>
<intersection>-87 1</intersection>
<intersection>-85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216.5,-87,228,-87</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>216.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>205.5,-85.5,216.5,-85.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>216.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216.5,-91.5,216.5,-89</points>
<intersection>-91.5 1</intersection>
<intersection>-89 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205.5,-91.5,216.5,-91.5</points>
<connection>
<GID>177</GID>
<name>OUT</name></connection>
<intersection>216.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216.5,-89,228,-89</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>216.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>208.5,-55,217,-55</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>208.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>208.5,-62,208.5,-55</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>-55 1</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,-105,225.5,-98.5</points>
<intersection>-105 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225.5,-105,230.5,-105</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,-98.5,225.5,-98.5</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,-98.5,212,-98</points>
<intersection>-98.5 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209.5,-98,212,-98</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>212,-98.5,214.5,-98.5</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>212 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-102,213,-100.5</points>
<intersection>-102 2</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213,-100.5,214.5,-100.5</points>
<connection>
<GID>179</GID>
<name>IN_2</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>212,-102,213,-102</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-17.2616,161.149,1206.74,-443.851</PageViewport></page 2>
<page 3>
<PageViewport>-17.2616,161.149,1206.74,-443.851</PageViewport></page 3>
<page 4>
<PageViewport>-17.2616,161.149,1206.74,-443.851</PageViewport></page 4>
<page 5>
<PageViewport>-17.2616,161.149,1206.74,-443.851</PageViewport></page 5>
<page 6>
<PageViewport>-17.2616,161.149,1206.74,-443.851</PageViewport></page 6>
<page 7>
<PageViewport>-17.2616,161.149,1206.74,-443.851</PageViewport></page 7>
<page 8>
<PageViewport>-17.2616,161.149,1206.74,-443.851</PageViewport></page 8>
<page 9>
<PageViewport>-17.2616,161.149,1206.74,-443.851</PageViewport></page 9></circuit>